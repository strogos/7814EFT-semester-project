
* Spice subcircuit definition for ADDFHX1


*.BIPOLAR
.GLOBAL VDD VSS

.subckt ANTENNA / A
DD1 A VDD pdio area=6.84e-13 pj=3.34e-06 m=1
DD0 VSS A ndio area=4.32e-13 pj=2.64e-06 m=1
.ends ANTENNA

.subckt ADDFHX1 CO S / A B CI
mn0 n0 A VSS VSS nmos1v w=0.34u l=0.1u
mn1 n0 B COb VSS nmos1v w=0.34u l=0.1u
mn10 n6 B n7 VSS nmos1v w=0.34u l=0.1u
mn11 n7 CI Sb VSS nmos1v w=0.34u l=0.1u
mn12 CO COb VSS VSS nmos1v w=0.43u l=0.1u
mn13 S Sb VSS VSS nmos1v w=0.43u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.34u l=0.1u
mn3 n2 B VSS VSS nmos1v w=0.34u l=0.1u
mn4 n2 CI COb VSS nmos1v w=0.34u l=0.1u
mn5 n4 A VSS VSS nmos1v w=0.34u l=0.1u
mn6 n4 B VSS VSS nmos1v w=0.34u l=0.1u
mn7 n4 CI VSS VSS nmos1v w=0.34u l=0.1u
mn8 n4 COb Sb VSS nmos1v w=0.34u l=0.1u
mn9 n6 A VSS VSS nmos1v w=0.34u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.52u l=0.1u
mp1 n1 B COb VDD pmos1v w=0.52u l=0.1u
mp10 n8 B n9 VDD pmos1v w=0.52u l=0.1u
mp11 n9 CI Sb VDD pmos1v w=0.52u l=0.1u
mp12 CO COb VDD VDD pmos1v w=0.65u l=0.1u
mp13 S Sb VDD VDD pmos1v w=0.65u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.52u l=0.1u
mp3 n3 B VDD VDD pmos1v w=0.52u l=0.1u
mp4 n3 CI COb VDD pmos1v w=0.52u l=0.1u
mp5 n5 A VDD VDD pmos1v w=0.52u l=0.1u
mp6 n5 B VDD VDD pmos1v w=0.52u l=0.1u
mp7 n5 CI VDD VDD pmos1v w=0.52u l=0.1u
mp8 n5 COb Sb VDD pmos1v w=0.52u l=0.1u
mp9 n8 A VDD VDD pmos1v w=0.52u l=0.1u
.ends ADDFHX1

* Spice subcircuit definition for ADDFHX2




.subckt ADDFHX2 CO S / A B CI
mn0 n0 A VSS VSS nmos1v w=0.34u l=0.1u
mn1 n0 B COb VSS nmos1v w=0.34u l=0.1u
mn10 n6 B n7 VSS nmos1v w=0.34u l=0.1u
mn11 n7 CI Sb VSS nmos1v w=0.34u l=0.1u
mn12 CO COb VSS VSS nmos1v w=0.86u l=0.1u
mn13 S Sb VSS VSS nmos1v w=0.86u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.34u l=0.1u
mn3 n2 B VSS VSS nmos1v w=0.34u l=0.1u
mn4 n2 CI COb VSS nmos1v w=0.34u l=0.1u
mn5 n4 A VSS VSS nmos1v w=0.34u l=0.1u
mn6 n4 B VSS VSS nmos1v w=0.34u l=0.1u
mn7 n4 CI VSS VSS nmos1v w=0.34u l=0.1u
mn8 n4 COb Sb VSS nmos1v w=0.34u l=0.1u
mn9 n6 A VSS VSS nmos1v w=0.34u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.52u l=0.1u
mp1 n1 B COb VDD pmos1v w=0.52u l=0.1u
mp10 n8 B n9 VDD pmos1v w=0.52u l=0.1u
mp11 n9 CI Sb VDD pmos1v w=0.52u l=0.1u
mp12 CO COb VDD VDD pmos1v w=1.3u l=0.1u
mp13 S Sb VDD VDD pmos1v w=1.3u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.52u l=0.1u
mp3 n3 B VDD VDD pmos1v w=0.52u l=0.1u
mp4 n3 CI COb VDD pmos1v w=0.52u l=0.1u
mp5 n5 A VDD VDD pmos1v w=0.52u l=0.1u
mp6 n5 B VDD VDD pmos1v w=0.52u l=0.1u
mp7 n5 CI VDD VDD pmos1v w=0.52u l=0.1u
mp8 n5 COb Sb VDD pmos1v w=0.52u l=0.1u
mp9 n8 A VDD VDD pmos1v w=0.52u l=0.1u
.ends ADDFHX2

* Spice subcircuit definition for ADDFHX4




.subckt ADDFHX4 CO S / A B CI
mn0 n0 A VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 B COb VSS nmos1v w=0.43u l=0.1u
mn10 n6 B n7 VSS nmos1v w=0.43u l=0.1u
mn11 n7 CI Sb VSS nmos1v w=0.43u l=0.1u
mn12 CO COb VSS VSS nmos1v w=1.72u l=0.1u
mn13 S Sb VSS VSS nmos1v w=1.72u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.43u l=0.1u
mn3 n2 B VSS VSS nmos1v w=0.43u l=0.1u
mn4 n2 CI COb VSS nmos1v w=0.43u l=0.1u
mn5 n4 A VSS VSS nmos1v w=0.43u l=0.1u
mn6 n4 B VSS VSS nmos1v w=0.43u l=0.1u
mn7 n4 CI VSS VSS nmos1v w=0.43u l=0.1u
mn8 n4 COb Sb VSS nmos1v w=0.43u l=0.1u
mn9 n6 A VSS VSS nmos1v w=0.43u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 B COb VDD pmos1v w=0.65u l=0.1u
mp10 n8 B n9 VDD pmos1v w=0.65u l=0.1u
mp11 n9 CI Sb VDD pmos1v w=0.65u l=0.1u
mp12 CO COb VDD VDD pmos1v w=2.6u l=0.1u
mp13 S Sb VDD VDD pmos1v w=2.6u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.65u l=0.1u
mp3 n3 B VDD VDD pmos1v w=0.65u l=0.1u
mp4 n3 CI COb VDD pmos1v w=0.65u l=0.1u
mp5 n5 A VDD VDD pmos1v w=0.65u l=0.1u
mp6 n5 B VDD VDD pmos1v w=0.65u l=0.1u
mp7 n5 CI VDD VDD pmos1v w=0.65u l=0.1u
mp8 n5 COb Sb VDD pmos1v w=0.65u l=0.1u
mp9 n8 A VDD VDD pmos1v w=0.65u l=0.1u
.ends ADDFHX4

* Spice subcircuit definition for ADDFHXL




.subckt ADDFHXL CO S / A B CI
mn0 n0 A VSS VSS nmos1v w=0.34u l=0.1u
mn1 n0 B COb VSS nmos1v w=0.34u l=0.1u
mn10 n6 B n7 VSS nmos1v w=0.34u l=0.1u
mn11 n7 CI Sb VSS nmos1v w=0.34u l=0.1u
mn12 CO COb VSS VSS nmos1v w=0.34u l=0.1u
mn13 S Sb VSS VSS nmos1v w=0.34u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.34u l=0.1u
mn3 n2 B VSS VSS nmos1v w=0.34u l=0.1u
mn4 n2 CI COb VSS nmos1v w=0.34u l=0.1u
mn5 n4 A VSS VSS nmos1v w=0.34u l=0.1u
mn6 n4 B VSS VSS nmos1v w=0.34u l=0.1u
mn7 n4 CI VSS VSS nmos1v w=0.34u l=0.1u
mn8 n4 COb Sb VSS nmos1v w=0.34u l=0.1u
mn9 n6 A VSS VSS nmos1v w=0.34u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.52u l=0.1u
mp1 n1 B COb VDD pmos1v w=0.52u l=0.1u
mp10 n8 B n9 VDD pmos1v w=0.52u l=0.1u
mp11 n9 CI Sb VDD pmos1v w=0.52u l=0.1u
mp12 CO COb VDD VDD pmos1v w=0.52u l=0.1u
mp13 S Sb VDD VDD pmos1v w=0.52u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.52u l=0.1u
mp3 n3 B VDD VDD pmos1v w=0.52u l=0.1u
mp4 n3 CI COb VDD pmos1v w=0.52u l=0.1u
mp5 n5 A VDD VDD pmos1v w=0.52u l=0.1u
mp6 n5 B VDD VDD pmos1v w=0.52u l=0.1u
mp7 n5 CI VDD VDD pmos1v w=0.52u l=0.1u
mp8 n5 COb Sb VDD pmos1v w=0.52u l=0.1u
mp9 n8 A VDD VDD pmos1v w=0.52u l=0.1u
.ends ADDFHXL

* Spice subcircuit definition for ADDFX1




.subckt ADDFX1 CO S / A B CI
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 B COb VSS nmos1v w=0.24u l=0.1u
mn10 n6 B n7 VSS nmos1v w=0.24u l=0.1u
mn11 n7 CI Sb VSS nmos1v w=0.24u l=0.1u
mn12 CO COb VSS VSS nmos1v w=0.43u l=0.1u
mn13 S Sb VSS VSS nmos1v w=0.43u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 B VSS VSS nmos1v w=0.24u l=0.1u
mn4 n2 CI COb VSS nmos1v w=0.24u l=0.1u
mn5 n4 A VSS VSS nmos1v w=0.24u l=0.1u
mn6 n4 B VSS VSS nmos1v w=0.24u l=0.1u
mn7 n4 CI VSS VSS nmos1v w=0.24u l=0.1u
mn8 n4 COb Sb VSS nmos1v w=0.24u l=0.1u
mn9 n6 A VSS VSS nmos1v w=0.24u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B COb VDD pmos1v w=0.36u l=0.1u
mp10 n8 B n9 VDD pmos1v w=0.36u l=0.1u
mp11 n9 CI Sb VDD pmos1v w=0.36u l=0.1u
mp12 CO COb VDD VDD pmos1v w=0.65u l=0.1u
mp13 S Sb VDD VDD pmos1v w=0.65u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 B VDD VDD pmos1v w=0.36u l=0.1u
mp4 n3 CI COb VDD pmos1v w=0.36u l=0.1u
mp5 n5 A VDD VDD pmos1v w=0.36u l=0.1u
mp6 n5 B VDD VDD pmos1v w=0.36u l=0.1u
mp7 n5 CI VDD VDD pmos1v w=0.36u l=0.1u
mp8 n5 COb Sb VDD pmos1v w=0.36u l=0.1u
mp9 n8 A VDD VDD pmos1v w=0.36u l=0.1u
.ends ADDFX1

* Spice subcircuit definition for ADDFX2




.subckt ADDFX2 CO S / A B CI
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 B COb VSS nmos1v w=0.24u l=0.1u
mn10 n6 B n7 VSS nmos1v w=0.24u l=0.1u
mn11 n7 CI Sb VSS nmos1v w=0.24u l=0.1u
mn12 CO COb VSS VSS nmos1v w=0.86u l=0.1u
mn13 S Sb VSS VSS nmos1v w=0.86u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 B VSS VSS nmos1v w=0.24u l=0.1u
mn4 n2 CI COb VSS nmos1v w=0.24u l=0.1u
mn5 n4 A VSS VSS nmos1v w=0.24u l=0.1u
mn6 n4 B VSS VSS nmos1v w=0.24u l=0.1u
mn7 n4 CI VSS VSS nmos1v w=0.24u l=0.1u
mn8 n4 COb Sb VSS nmos1v w=0.24u l=0.1u
mn9 n6 A VSS VSS nmos1v w=0.24u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B COb VDD pmos1v w=0.36u l=0.1u
mp10 n8 B n9 VDD pmos1v w=0.36u l=0.1u
mp11 n9 CI Sb VDD pmos1v w=0.36u l=0.1u
mp12 CO COb VDD VDD pmos1v w=1.3u l=0.1u
mp13 S Sb VDD VDD pmos1v w=1.3u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 B VDD VDD pmos1v w=0.36u l=0.1u
mp4 n3 CI COb VDD pmos1v w=0.36u l=0.1u
mp5 n5 A VDD VDD pmos1v w=0.36u l=0.1u
mp6 n5 B VDD VDD pmos1v w=0.36u l=0.1u
mp7 n5 CI VDD VDD pmos1v w=0.36u l=0.1u
mp8 n5 COb Sb VDD pmos1v w=0.36u l=0.1u
mp9 n8 A VDD VDD pmos1v w=0.36u l=0.1u
.ends ADDFX2

* Spice subcircuit definition for ADDFX4




.subckt ADDFX4 CO S / A B CI
mn0 n0 A VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 B COb VSS nmos1v w=0.43u l=0.1u
mn10 n6 B n7 VSS nmos1v w=0.43u l=0.1u
mn11 n7 CI Sb VSS nmos1v w=0.43u l=0.1u
mn12 CO COb VSS VSS nmos1v w=1.72u l=0.1u
mn13 S Sb VSS VSS nmos1v w=1.72u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.43u l=0.1u
mn3 n2 B VSS VSS nmos1v w=0.43u l=0.1u
mn4 n2 CI COb VSS nmos1v w=0.43u l=0.1u
mn5 n4 A VSS VSS nmos1v w=0.43u l=0.1u
mn6 n4 B VSS VSS nmos1v w=0.43u l=0.1u
mn7 n4 CI VSS VSS nmos1v w=0.43u l=0.1u
mn8 n4 COb Sb VSS nmos1v w=0.43u l=0.1u
mn9 n6 A VSS VSS nmos1v w=0.43u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 B COb VDD pmos1v w=0.65u l=0.1u
mp10 n8 B n9 VDD pmos1v w=0.65u l=0.1u
mp11 n9 CI Sb VDD pmos1v w=0.65u l=0.1u
mp12 CO COb VDD VDD pmos1v w=2.6u l=0.1u
mp13 S Sb VDD VDD pmos1v w=2.6u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.65u l=0.1u
mp3 n3 B VDD VDD pmos1v w=0.65u l=0.1u
mp4 n3 CI COb VDD pmos1v w=0.65u l=0.1u
mp5 n5 A VDD VDD pmos1v w=0.65u l=0.1u
mp6 n5 B VDD VDD pmos1v w=0.65u l=0.1u
mp7 n5 CI VDD VDD pmos1v w=0.65u l=0.1u
mp8 n5 COb Sb VDD pmos1v w=0.65u l=0.1u
mp9 n8 A VDD VDD pmos1v w=0.65u l=0.1u
.ends ADDFX4

* Spice subcircuit definition for ADDFXL




.subckt ADDFXL CO S / A B CI
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 B COb VSS nmos1v w=0.24u l=0.1u
mn10 n6 B n7 VSS nmos1v w=0.24u l=0.1u
mn11 n7 CI Sb VSS nmos1v w=0.24u l=0.1u
mn12 CO COb VSS VSS nmos1v w=0.24u l=0.1u
mn13 S Sb VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 B VSS VSS nmos1v w=0.24u l=0.1u
mn4 n2 CI COb VSS nmos1v w=0.24u l=0.1u
mn5 n4 A VSS VSS nmos1v w=0.24u l=0.1u
mn6 n4 B VSS VSS nmos1v w=0.24u l=0.1u
mn7 n4 CI VSS VSS nmos1v w=0.24u l=0.1u
mn8 n4 COb Sb VSS nmos1v w=0.24u l=0.1u
mn9 n6 A VSS VSS nmos1v w=0.24u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B COb VDD pmos1v w=0.36u l=0.1u
mp10 n8 B n9 VDD pmos1v w=0.36u l=0.1u
mp11 n9 CI Sb VDD pmos1v w=0.36u l=0.1u
mp12 CO COb VDD VDD pmos1v w=0.36u l=0.1u
mp13 S Sb VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 B VDD VDD pmos1v w=0.36u l=0.1u
mp4 n3 CI COb VDD pmos1v w=0.36u l=0.1u
mp5 n5 A VDD VDD pmos1v w=0.36u l=0.1u
mp6 n5 B VDD VDD pmos1v w=0.36u l=0.1u
mp7 n5 CI VDD VDD pmos1v w=0.36u l=0.1u
mp8 n5 COb Sb VDD pmos1v w=0.36u l=0.1u
mp9 n8 A VDD VDD pmos1v w=0.36u l=0.1u
.ends ADDFXL

* Spice subcircuit definition for ADDHX1




.subckt ADDHX1 CO S / A B
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 B Sb VSS nmos1v w=0.24u l=0.1u
mn4 n0 n1 Sb VSS nmos1v w=0.24u l=0.1u
mn5 S Sb VSS VSS nmos1v w=0.43u l=0.1u
mn6 n4 A VSS VSS nmos1v w=0.24u l=0.1u
mn7 n4 B COb VSS nmos1v w=0.24u l=0.1u
mn8 CO COb VSS VSS nmos1v w=0.43u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 n1 Sb VDD pmos1v w=0.36u l=0.1u
mp4 n0 B Sb VDD pmos1v w=0.36u l=0.1u
mp5 S Sb VDD VDD pmos1v w=0.65u l=0.1u
mp6 COb A VDD VDD pmos1v w=0.36u l=0.1u
mp7 COb B VDD VDD pmos1v w=0.36u l=0.1u
mp8 CO COb VDD VDD pmos1v w=0.65u l=0.1u
.ends ADDHX1

* Spice subcircuit definition for ADDHX2




.subckt ADDHX2 CO S / A B
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 B Sb VSS nmos1v w=0.24u l=0.1u
mn4 n0 n1 Sb VSS nmos1v w=0.24u l=0.1u
mn5 S Sb VSS VSS nmos1v w=0.86u l=0.1u
mn6 n4 A VSS VSS nmos1v w=0.24u l=0.1u
mn7 n4 B COb VSS nmos1v w=0.24u l=0.1u
mn8 CO COb VSS VSS nmos1v w=0.86u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 n1 Sb VDD pmos1v w=0.36u l=0.1u
mp4 n0 B Sb VDD pmos1v w=0.36u l=0.1u
mp5 S Sb VDD VDD pmos1v w=1.3u l=0.1u
mp6 COb A VDD VDD pmos1v w=0.36u l=0.1u
mp7 COb B VDD VDD pmos1v w=0.36u l=0.1u
mp8 CO COb VDD VDD pmos1v w=1.3u l=0.1u
.ends ADDHX2

* Spice subcircuit definition for ADDHX4




.subckt ADDHX4 CO S / A B
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=0.43u l=0.1u
mn3 n2 B Sb VSS nmos1v w=0.43u l=0.1u
mn4 n0 n1 Sb VSS nmos1v w=0.43u l=0.1u
mn5 S Sb VSS VSS nmos1v w=1.72u l=0.1u
mn6 n4 A VSS VSS nmos1v w=0.43u l=0.1u
mn7 n4 B COb VSS nmos1v w=0.43u l=0.1u
mn8 CO COb VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 n0 VDD VDD pmos1v w=0.65u l=0.1u
mp3 n3 n1 Sb VDD pmos1v w=0.65u l=0.1u
mp4 n0 B Sb VDD pmos1v w=0.65u l=0.1u
mp5 S Sb VDD VDD pmos1v w=2.6u l=0.1u
mp6 COb A VDD VDD pmos1v w=0.65u l=0.1u
mp7 COb B VDD VDD pmos1v w=0.65u l=0.1u
mp8 CO COb VDD VDD pmos1v w=2.6u l=0.1u
.ends ADDHX4

* Spice subcircuit definition for ADDHXL




.subckt ADDHXL CO S / A B
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 B Sb VSS nmos1v w=0.24u l=0.1u
mn4 n0 n1 Sb VSS nmos1v w=0.24u l=0.1u
mn5 S Sb VSS VSS nmos1v w=0.24u l=0.1u
mn6 n4 A VSS VSS nmos1v w=0.24u l=0.1u
mn7 n4 B COb VSS nmos1v w=0.24u l=0.1u
mn8 CO COb VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 n1 Sb VDD pmos1v w=0.36u l=0.1u
mp4 n0 B Sb VDD pmos1v w=0.36u l=0.1u
mp5 S Sb VDD VDD pmos1v w=0.36u l=0.1u
mp6 COb A VDD VDD pmos1v w=0.36u l=0.1u
mp7 COb B VDD VDD pmos1v w=0.36u l=0.1u
mp8 CO COb VDD VDD pmos1v w=0.36u l=0.1u
.ends ADDHXL

* Spice subcircuit definition for AND2X1




.subckt AND2X1 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 B n0 VSS nmos1v w=0.24u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends AND2X1

* Spice subcircuit definition for AND2X2




.subckt AND2X2 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 B n0 VSS nmos1v w=0.24u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends AND2X2

* Spice subcircuit definition for AND2X4




.subckt AND2X4 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.43u l=0.1u
mn1 n1 B n0 VSS nmos1v w=0.43u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 n0 B VDD VDD pmos1v w=0.65u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends AND2X4

* Spice subcircuit definition for AND2X6




.subckt AND2X6 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n1 B n0 VSS nmos1v w=0.86u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=2.58u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n0 B VDD VDD pmos1v w=1.3u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=3.9u l=0.1u
.ends AND2X6

* Spice subcircuit definition for AND2X8




.subckt AND2X8 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n1 B n0 VSS nmos1v w=0.86u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=3.44u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n0 B VDD VDD pmos1v w=1.3u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=5.2u l=0.1u
.ends AND2X8

* Spice subcircuit definition for AND2XL




.subckt AND2XL Y / A B
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 B n0 VSS nmos1v w=0.24u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
.ends AND2XL

* Spice subcircuit definition for AND3X1




.subckt AND3X1 Y / A B C
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 B n2 VSS nmos1v w=0.24u l=0.1u
mn2 n2 C n0 VSS nmos1v w=0.24u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n0 C VDD VDD pmos1v w=0.36u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends AND3X1

* Spice subcircuit definition for AND3X2




.subckt AND3X2 Y / A B C
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 B n2 VSS nmos1v w=0.24u l=0.1u
mn2 n2 C n0 VSS nmos1v w=0.24u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n0 C VDD VDD pmos1v w=0.36u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends AND3X2

* Spice subcircuit definition for AND3X4




.subckt AND3X4 Y / A B C
mn0 n1 A VSS VSS nmos1v w=0.43u l=0.1u
mn1 n1 B n2 VSS nmos1v w=0.43u l=0.1u
mn2 n2 C n0 VSS nmos1v w=0.43u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 n0 B VDD VDD pmos1v w=0.65u l=0.1u
mp2 n0 C VDD VDD pmos1v w=0.65u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends AND3X4

* Spice subcircuit definition for AND3X6




.subckt AND3X6 Y / A B C
mn0 n1 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n1 B n2 VSS nmos1v w=0.86u l=0.1u
mn2 n2 C n0 VSS nmos1v w=0.86u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=2.58u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n0 B VDD VDD pmos1v w=1.3u l=0.1u
mp2 n0 C VDD VDD pmos1v w=1.3u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=3.9u l=0.1u
.ends AND3X6

* Spice subcircuit definition for AND3X8




.subckt AND3X8 Y / A B C
mn0 n1 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n1 B n2 VSS nmos1v w=0.86u l=0.1u
mn2 n2 C n0 VSS nmos1v w=0.86u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=3.44u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n0 B VDD VDD pmos1v w=1.3u l=0.1u
mp2 n0 C VDD VDD pmos1v w=1.3u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=5.2u l=0.1u
.ends AND3X8

* Spice subcircuit definition for AND3XL




.subckt AND3XL Y / A B C
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 B n2 VSS nmos1v w=0.24u l=0.1u
mn2 n2 C n0 VSS nmos1v w=0.24u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n0 C VDD VDD pmos1v w=0.36u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
.ends AND3XL

* Spice subcircuit definition for AND4X1




.subckt AND4X1 Y / A B C D
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 B n2 VSS nmos1v w=0.24u l=0.1u
mn2 n2 C n3 VSS nmos1v w=0.24u l=0.1u
mn3 n3 D n0 VSS nmos1v w=0.24u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n0 C VDD VDD pmos1v w=0.36u l=0.1u
mp3 n0 D VDD VDD pmos1v w=0.36u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends AND4X1

* Spice subcircuit definition for AND4X2




.subckt AND4X2 Y / A B C D
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 B n2 VSS nmos1v w=0.24u l=0.1u
mn2 n2 C n3 VSS nmos1v w=0.24u l=0.1u
mn3 n3 D n0 VSS nmos1v w=0.24u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n0 C VDD VDD pmos1v w=0.36u l=0.1u
mp3 n0 D VDD VDD pmos1v w=0.36u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends AND4X2

* Spice subcircuit definition for AND4X4




.subckt AND4X4 Y / A B C D
mn0 n1 A VSS VSS nmos1v w=0.43u l=0.1u
mn1 n1 B n2 VSS nmos1v w=0.43u l=0.1u
mn2 n2 C n3 VSS nmos1v w=0.43u l=0.1u
mn3 n3 D n0 VSS nmos1v w=0.43u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 n0 B VDD VDD pmos1v w=0.65u l=0.1u
mp2 n0 C VDD VDD pmos1v w=0.65u l=0.1u
mp3 n0 D VDD VDD pmos1v w=0.65u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends AND4X4

* Spice subcircuit definition for AND4X6




.subckt AND4X6 Y / A B C D
mn0 n1 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n1 B n2 VSS nmos1v w=0.86u l=0.1u
mn2 n2 C n3 VSS nmos1v w=0.86u l=0.1u
mn3 n3 D n0 VSS nmos1v w=0.86u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=2.58u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n0 B VDD VDD pmos1v w=1.3u l=0.1u
mp2 n0 C VDD VDD pmos1v w=1.3u l=0.1u
mp3 n0 D VDD VDD pmos1v w=1.3u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=3.9u l=0.1u
.ends AND4X6

* Spice subcircuit definition for AND4X8




.subckt AND4X8 Y / A B C D
mn0 n1 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n1 B n2 VSS nmos1v w=0.86u l=0.1u
mn2 n2 C n3 VSS nmos1v w=0.86u l=0.1u
mn3 n3 D n0 VSS nmos1v w=0.86u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=3.44u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n0 B VDD VDD pmos1v w=1.3u l=0.1u
mp2 n0 C VDD VDD pmos1v w=1.3u l=0.1u
mp3 n0 D VDD VDD pmos1v w=1.3u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=5.2u l=0.1u
.ends AND4X8

* Spice subcircuit definition for AND4XL




.subckt AND4XL Y / A B C D
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 B n2 VSS nmos1v w=0.24u l=0.1u
mn2 n2 C n3 VSS nmos1v w=0.24u l=0.1u
mn3 n3 D n0 VSS nmos1v w=0.24u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n0 C VDD VDD pmos1v w=0.36u l=0.1u
mp3 n0 D VDD VDD pmos1v w=0.36u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
.ends AND4XL

* Spice subcircuit definition for AO21X1




.subckt AO21X1 Y / A0 A1 B0
mn0 n1 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1 n0 VSS nmos1v w=0.24u l=0.1u
mn2 n0 B0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n2 B0 n0 VDD pmos1v w=0.36u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends AO21X1

* Spice subcircuit definition for AO21X2




.subckt AO21X2 Y / A0 A1 B0
mn0 n1 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1 n0 VSS nmos1v w=0.24u l=0.1u
mn2 n0 B0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n2 B0 n0 VDD pmos1v w=0.36u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends AO21X2

* Spice subcircuit definition for AO21X4




.subckt AO21X4 Y / A0 A1 B0
mn0 n1 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n1 A1 n0 VSS nmos1v w=0.43u l=0.1u
mn2 n0 B0 VSS VSS nmos1v w=0.43u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n2 B0 n0 VDD pmos1v w=0.65u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends AO21X4

* Spice subcircuit definition for AO21XL




.subckt AO21XL Y / A0 A1 B0
mn0 n1 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1 n0 VSS nmos1v w=0.24u l=0.1u
mn2 n0 B0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n2 B0 n0 VDD pmos1v w=0.36u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
.ends AO21XL

* Spice subcircuit definition for AO22X1




.subckt AO22X1 Y / A0 A1 B0 B1
mn0 n1 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1 n0 VSS nmos1v w=0.24u l=0.1u
mn2 n2 B0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 B1 n0 VSS nmos1v w=0.24u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n3 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n3 A1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 B0 n0 VDD pmos1v w=0.36u l=0.1u
mp3 n3 B1 n0 VDD pmos1v w=0.36u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends AO22X1

* Spice subcircuit definition for AO22X2




.subckt AO22X2 Y / A0 A1 B0 B1
mn0 n1 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1 n0 VSS nmos1v w=0.24u l=0.1u
mn2 n2 B0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 B1 n0 VSS nmos1v w=0.24u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n3 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n3 A1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 B0 n0 VDD pmos1v w=0.36u l=0.1u
mp3 n3 B1 n0 VDD pmos1v w=0.36u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends AO22X2

* Spice subcircuit definition for AO22X4




.subckt AO22X4 Y / A0 A1 B0 B1
mn0 n1 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n1 A1 n0 VSS nmos1v w=0.43u l=0.1u
mn2 n2 B0 VSS VSS nmos1v w=0.43u l=0.1u
mn3 n2 B1 n0 VSS nmos1v w=0.43u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n3 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n3 A1 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n3 B0 n0 VDD pmos1v w=0.65u l=0.1u
mp3 n3 B1 n0 VDD pmos1v w=0.65u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends AO22X4

* Spice subcircuit definition for AO22XL




.subckt AO22XL Y / A0 A1 B0 B1
mn0 n1 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1 n0 VSS nmos1v w=0.24u l=0.1u
mn2 n2 B0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 B1 n0 VSS nmos1v w=0.24u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n3 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n3 A1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 B0 n0 VDD pmos1v w=0.36u l=0.1u
mp3 n3 B1 n0 VDD pmos1v w=0.36u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
.ends AO22XL

* Spice subcircuit definition for AOI211X1




.subckt AOI211X1 Y / A0 A1 B0 C0
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=0.43u l=0.1u
mn2 Y B0 VSS VSS nmos1v w=0.43u l=0.1u
mn3 Y C0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 A1 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n1 B0 n2 VDD pmos1v w=0.65u l=0.1u
mp3 n2 C0 Y VDD pmos1v w=0.65u l=0.1u
.ends AOI211X1

* Spice subcircuit definition for AOI211X2




.subckt AOI211X2 Y / A0 A1 B0 C0
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=0.86u l=0.1u
mn2 Y B0 VSS VSS nmos1v w=0.86u l=0.1u
mn3 Y C0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n1 A1 VDD VDD pmos1v w=1.3u l=0.1u
mp2 n1 B0 n2 VDD pmos1v w=1.3u l=0.1u
mp3 n2 C0 Y VDD pmos1v w=1.3u l=0.1u
.ends AOI211X2

* Spice subcircuit definition for AOI211X4




.subckt AOI211X4 Y / A0 A1 B0 C0
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=1.72u l=0.1u
mn2 Y B0 VSS VSS nmos1v w=1.72u l=0.1u
mn3 Y C0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n1 A1 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n1 B0 n2 VDD pmos1v w=2.6u l=0.1u
mp3 n2 C0 Y VDD pmos1v w=2.6u l=0.1u
.ends AOI211X4

* Spice subcircuit definition for AOI211XL




.subckt AOI211XL Y / A0 A1 B0 C0
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=0.24u l=0.1u
mn2 Y B0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 Y C0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n1 B0 n2 VDD pmos1v w=0.36u l=0.1u
mp3 n2 C0 Y VDD pmos1v w=0.36u l=0.1u
.ends AOI211XL

* Spice subcircuit definition for AOI21X1




.subckt AOI21X1 Y / A0 A1 B0
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=0.43u l=0.1u
mn2 Y B0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 A1 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n1 B0 Y VDD pmos1v w=0.65u l=0.1u
.ends AOI21X1

* Spice subcircuit definition for AOI21X2




.subckt AOI21X2 Y / A0 A1 B0
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=0.86u l=0.1u
mn2 Y B0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n1 A1 VDD VDD pmos1v w=1.3u l=0.1u
mp2 n1 B0 Y VDD pmos1v w=1.3u l=0.1u
.ends AOI21X2

* Spice subcircuit definition for AOI21X4




.subckt AOI21X4 Y / A0 A1 B0
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=1.72u l=0.1u
mn2 Y B0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n1 A1 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n1 B0 Y VDD pmos1v w=2.6u l=0.1u
.ends AOI21X4

* Spice subcircuit definition for AOI21XL




.subckt AOI21XL Y / A0 A1 B0
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=0.24u l=0.1u
mn2 Y B0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n1 B0 Y VDD pmos1v w=0.36u l=0.1u
.ends AOI21XL

* Spice subcircuit definition for AOI221X1




.subckt AOI221X1 Y / A0 A1 B0 B1 C0
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=0.43u l=0.1u
mn2 n1 B0 VSS VSS nmos1v w=0.43u l=0.1u
mn3 n1 B1 Y VSS nmos1v w=0.43u l=0.1u
mn4 Y C0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n2 B0 n3 VDD pmos1v w=0.65u l=0.1u
mp3 n2 B1 n3 VDD pmos1v w=0.65u l=0.1u
mp4 n3 C0 Y VDD pmos1v w=0.65u l=0.1u
.ends AOI221X1

* Spice subcircuit definition for AOI221X2




.subckt AOI221X2 Y / A0 A1 B0 B1 C0
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=0.86u l=0.1u
mn2 n1 B0 VSS VSS nmos1v w=0.86u l=0.1u
mn3 n1 B1 Y VSS nmos1v w=0.86u l=0.1u
mn4 Y C0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=1.3u l=0.1u
mp2 n2 B0 n3 VDD pmos1v w=1.3u l=0.1u
mp3 n2 B1 n3 VDD pmos1v w=1.3u l=0.1u
mp4 n3 C0 Y VDD pmos1v w=1.3u l=0.1u
.ends AOI221X2

* Spice subcircuit definition for AOI221X4




.subckt AOI221X4 Y / A0 A1 B0 B1 C0
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=1.72u l=0.1u
mn2 n1 B0 VSS VSS nmos1v w=1.72u l=0.1u
mn3 n1 B1 Y VSS nmos1v w=1.72u l=0.1u
mn4 Y C0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n2 B0 n3 VDD pmos1v w=2.6u l=0.1u
mp3 n2 B1 n3 VDD pmos1v w=2.6u l=0.1u
mp4 n3 C0 Y VDD pmos1v w=2.6u l=0.1u
.ends AOI221X4

* Spice subcircuit definition for AOI221XL




.subckt AOI221XL Y / A0 A1 B0 B1 C0
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=0.24u l=0.1u
mn2 n1 B0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n1 B1 Y VSS nmos1v w=0.24u l=0.1u
mn4 Y C0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n2 B0 n3 VDD pmos1v w=0.36u l=0.1u
mp3 n2 B1 n3 VDD pmos1v w=0.36u l=0.1u
mp4 n3 C0 Y VDD pmos1v w=0.36u l=0.1u
.ends AOI221XL

* Spice subcircuit definition for AOI222X1




.subckt AOI222X1 Y / A0 A1 B0 B1 C0 C1
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=0.43u l=0.1u
mn2 n1 B0 VSS VSS nmos1v w=0.43u l=0.1u
mn3 n1 B1 Y VSS nmos1v w=0.43u l=0.1u
mn4 n2 C0 VSS VSS nmos1v w=0.43u l=0.1u
mn5 n2 C1 Y VSS nmos1v w=0.43u l=0.1u
mp0 n3 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n3 A1 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n3 B0 n4 VDD pmos1v w=0.65u l=0.1u
mp3 n3 B1 n4 VDD pmos1v w=0.65u l=0.1u
mp4 n4 C0 Y VDD pmos1v w=0.65u l=0.1u
mp5 n4 C1 Y VDD pmos1v w=0.65u l=0.1u
.ends AOI222X1

* Spice subcircuit definition for AOI222X2




.subckt AOI222X2 Y / A0 A1 B0 B1 C0 C1
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=0.86u l=0.1u
mn2 n1 B0 VSS VSS nmos1v w=0.86u l=0.1u
mn3 n1 B1 Y VSS nmos1v w=0.86u l=0.1u
mn4 n2 C0 VSS VSS nmos1v w=0.86u l=0.1u
mn5 n2 C1 Y VSS nmos1v w=0.86u l=0.1u
mp0 n3 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n3 A1 VDD VDD pmos1v w=1.3u l=0.1u
mp2 n3 B0 n4 VDD pmos1v w=1.3u l=0.1u
mp3 n3 B1 n4 VDD pmos1v w=1.3u l=0.1u
mp4 n4 C0 Y VDD pmos1v w=1.3u l=0.1u
mp5 n4 C1 Y VDD pmos1v w=1.3u l=0.1u
.ends AOI222X2

* Spice subcircuit definition for AOI222X4




.subckt AOI222X4 Y / A0 A1 B0 B1 C0 C1
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=1.72u l=0.1u
mn2 n1 B0 VSS VSS nmos1v w=1.72u l=0.1u
mn3 n1 B1 Y VSS nmos1v w=1.72u l=0.1u
mn4 n2 C0 VSS VSS nmos1v w=1.72u l=0.1u
mn5 n2 C1 Y VSS nmos1v w=1.72u l=0.1u
mp0 n3 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n3 A1 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n3 B0 n4 VDD pmos1v w=2.6u l=0.1u
mp3 n3 B1 n4 VDD pmos1v w=2.6u l=0.1u
mp4 n4 C0 Y VDD pmos1v w=2.6u l=0.1u
mp5 n4 C1 Y VDD pmos1v w=2.6u l=0.1u
.ends AOI222X4

* Spice subcircuit definition for AOI222XL




.subckt AOI222XL Y / A0 A1 B0 B1 C0 C1
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=0.24u l=0.1u
mn2 n1 B0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n1 B1 Y VSS nmos1v w=0.24u l=0.1u
mn4 n2 C0 VSS VSS nmos1v w=0.24u l=0.1u
mn5 n2 C1 Y VSS nmos1v w=0.24u l=0.1u
mp0 n3 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n3 A1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 B0 n4 VDD pmos1v w=0.36u l=0.1u
mp3 n3 B1 n4 VDD pmos1v w=0.36u l=0.1u
mp4 n4 C0 Y VDD pmos1v w=0.36u l=0.1u
mp5 n4 C1 Y VDD pmos1v w=0.36u l=0.1u
.ends AOI222XL

* Spice subcircuit definition for AOI22X1




.subckt AOI22X1 Y / A0 A1 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=0.43u l=0.1u
mn2 n1 B0 VSS VSS nmos1v w=0.43u l=0.1u
mn3 n1 B1 Y VSS nmos1v w=0.43u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n2 B0 Y VDD pmos1v w=0.65u l=0.1u
mp3 n2 B1 Y VDD pmos1v w=0.65u l=0.1u
.ends AOI22X1

* Spice subcircuit definition for AOI22X2




.subckt AOI22X2 Y / A0 A1 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=0.86u l=0.1u
mn2 n1 B0 VSS VSS nmos1v w=0.86u l=0.1u
mn3 n1 B1 Y VSS nmos1v w=0.86u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=1.3u l=0.1u
mp2 n2 B0 Y VDD pmos1v w=1.3u l=0.1u
mp3 n2 B1 Y VDD pmos1v w=1.3u l=0.1u
.ends AOI22X2

* Spice subcircuit definition for AOI22X4




.subckt AOI22X4 Y / A0 A1 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=1.72u l=0.1u
mn2 n1 B0 VSS VSS nmos1v w=1.72u l=0.1u
mn3 n1 B1 Y VSS nmos1v w=1.72u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n2 B0 Y VDD pmos1v w=2.6u l=0.1u
mp3 n2 B1 Y VDD pmos1v w=2.6u l=0.1u
.ends AOI22X4

* Spice subcircuit definition for AOI22XL




.subckt AOI22XL Y / A0 A1 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 Y VSS nmos1v w=0.24u l=0.1u
mn2 n1 B0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n1 B1 Y VSS nmos1v w=0.24u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n2 B0 Y VDD pmos1v w=0.36u l=0.1u
mp3 n2 B1 Y VDD pmos1v w=0.36u l=0.1u
.ends AOI22XL

* Spice subcircuit definition for AOI2BB1X1




.subckt AOI2BB1X1 Y / A0N A1N B0
mn0 n0 A0N VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1N VSS VSS nmos1v w=0.24u l=0.1u
mn2 Y B0 VSS VSS nmos1v w=0.43u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n1 A0N VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1N n0 VDD pmos1v w=0.36u l=0.1u
mp2 n2 B0 VDD VDD pmos1v w=0.65u l=0.1u
mp3 n2 n0 Y VDD pmos1v w=0.65u l=0.1u
.ends AOI2BB1X1

* Spice subcircuit definition for AOI2BB1X2




.subckt AOI2BB1X2 Y / A0N A1N B0
mn0 n0 A0N VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1N VSS VSS nmos1v w=0.24u l=0.1u
mn2 Y B0 VSS VSS nmos1v w=0.86u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n1 A0N VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1N n0 VDD pmos1v w=0.36u l=0.1u
mp2 n2 B0 VDD VDD pmos1v w=1.3u l=0.1u
mp3 n2 n0 Y VDD pmos1v w=1.3u l=0.1u
.ends AOI2BB1X2

* Spice subcircuit definition for AOI2BB1X4




.subckt AOI2BB1X4 Y / A0N A1N B0
mn0 n0 A0N VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1N VSS VSS nmos1v w=0.43u l=0.1u
mn2 Y B0 VSS VSS nmos1v w=1.72u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n1 A0N VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 A1N n0 VDD pmos1v w=0.65u l=0.1u
mp2 n2 B0 VDD VDD pmos1v w=2.6u l=0.1u
mp3 n2 n0 Y VDD pmos1v w=2.6u l=0.1u
.ends AOI2BB1X4

* Spice subcircuit definition for AOI2BB1XL




.subckt AOI2BB1XL Y / A0N A1N B0
mn0 n0 A0N VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1N VSS VSS nmos1v w=0.24u l=0.1u
mn2 Y B0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n1 A0N VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1N n0 VDD pmos1v w=0.36u l=0.1u
mp2 n2 B0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n2 n0 Y VDD pmos1v w=0.36u l=0.1u
.ends AOI2BB1XL

* Spice subcircuit definition for AOI2BB2X1




.subckt AOI2BB2X1 Y / A0N A1N B0 B1
mn0 n0 A0N VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1N VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=0.43u l=0.1u
mn3 n2 n1 Y VSS nmos1v w=0.43u l=0.1u
mn4 n3 B0 VSS VSS nmos1v w=0.43u l=0.1u
mn5 n3 B1 Y VSS nmos1v w=0.43u l=0.1u
mp0 n0 A0N VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1N VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 n0 VDD VDD pmos1v w=0.65u l=0.1u
mp3 n4 n1 VDD VDD pmos1v w=0.65u l=0.1u
mp4 n4 B0 Y VDD pmos1v w=0.65u l=0.1u
mp5 n4 B1 Y VDD pmos1v w=0.65u l=0.1u
.ends AOI2BB2X1

* Spice subcircuit definition for AOI2BB2X2




.subckt AOI2BB2X2 Y / A0N A1N B0 B1
mn0 n0 A0N VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1N VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=0.86u l=0.1u
mn3 n2 n1 Y VSS nmos1v w=0.86u l=0.1u
mn4 n3 B0 VSS VSS nmos1v w=0.86u l=0.1u
mn5 n3 B1 Y VSS nmos1v w=0.86u l=0.1u
mp0 n0 A0N VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1N VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 n0 VDD VDD pmos1v w=1.3u l=0.1u
mp3 n4 n1 VDD VDD pmos1v w=1.3u l=0.1u
mp4 n4 B0 Y VDD pmos1v w=1.3u l=0.1u
mp5 n4 B1 Y VDD pmos1v w=1.3u l=0.1u
.ends AOI2BB2X2

* Spice subcircuit definition for AOI2BB2X4




.subckt AOI2BB2X4 Y / A0N A1N B0 B1
mn0 n0 A0N VSS VSS nmos1v w=0.43u l=0.1u
mn1 n1 A1N VSS VSS nmos1v w=0.43u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=1.72u l=0.1u
mn3 n2 n1 Y VSS nmos1v w=1.72u l=0.1u
mn4 n3 B0 VSS VSS nmos1v w=1.72u l=0.1u
mn5 n3 B1 Y VSS nmos1v w=1.72u l=0.1u
mp0 n0 A0N VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 A1N VDD VDD pmos1v w=0.65u l=0.1u
mp2 n4 n0 VDD VDD pmos1v w=2.6u l=0.1u
mp3 n4 n1 VDD VDD pmos1v w=2.6u l=0.1u
mp4 n4 B0 Y VDD pmos1v w=2.6u l=0.1u
mp5 n4 B1 Y VDD pmos1v w=2.6u l=0.1u
.ends AOI2BB2X4

* Spice subcircuit definition for AOI2BB2XL




.subckt AOI2BB2XL Y / A0N A1N B0 B1
mn0 n0 A0N VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1N VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 n1 Y VSS nmos1v w=0.24u l=0.1u
mn4 n3 B0 VSS VSS nmos1v w=0.24u l=0.1u
mn5 n3 B1 Y VSS nmos1v w=0.24u l=0.1u
mp0 n0 A0N VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1N VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp4 n4 B0 Y VDD pmos1v w=0.36u l=0.1u
mp5 n4 B1 Y VDD pmos1v w=0.36u l=0.1u
.ends AOI2BB2XL

* Spice subcircuit definition for AOI31X1




.subckt AOI31X1 Y / A0 A1 A2 B0
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 n1 VSS nmos1v w=0.43u l=0.1u
mn2 n1 A2 Y VSS nmos1v w=0.43u l=0.1u
mn3 Y B0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n2 A2 VDD VDD pmos1v w=0.65u l=0.1u
mp3 n2 B0 Y VDD pmos1v w=0.65u l=0.1u
.ends AOI31X1

* Spice subcircuit definition for AOI31X2




.subckt AOI31X2 Y / A0 A1 A2 B0
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 n1 VSS nmos1v w=0.86u l=0.1u
mn2 n1 A2 Y VSS nmos1v w=0.86u l=0.1u
mn3 Y B0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=1.3u l=0.1u
mp2 n2 A2 VDD VDD pmos1v w=1.3u l=0.1u
mp3 n2 B0 Y VDD pmos1v w=1.3u l=0.1u
.ends AOI31X2

* Spice subcircuit definition for AOI31X4




.subckt AOI31X4 Y / A0 A1 A2 B0
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 n1 VSS nmos1v w=1.72u l=0.1u
mn2 n1 A2 Y VSS nmos1v w=1.72u l=0.1u
mn3 Y B0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n2 A2 VDD VDD pmos1v w=2.6u l=0.1u
mp3 n2 B0 Y VDD pmos1v w=2.6u l=0.1u
.ends AOI31X4

* Spice subcircuit definition for AOI31XL




.subckt AOI31XL Y / A0 A1 A2 B0
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 n1 VSS nmos1v w=0.24u l=0.1u
mn2 n1 A2 Y VSS nmos1v w=0.24u l=0.1u
mn3 Y B0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 A1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n2 A2 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n2 B0 Y VDD pmos1v w=0.36u l=0.1u
.ends AOI31XL

* Spice subcircuit definition for AOI32X1




.subckt AOI32X1 Y / A0 A1 A2 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 n1 VSS nmos1v w=0.43u l=0.1u
mn2 n1 A2 Y VSS nmos1v w=0.43u l=0.1u
mn3 n2 B0 VSS VSS nmos1v w=0.43u l=0.1u
mn4 n2 B1 Y VSS nmos1v w=0.43u l=0.1u
mp0 n3 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n3 A1 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n3 A2 VDD VDD pmos1v w=0.65u l=0.1u
mp3 n3 B0 Y VDD pmos1v w=0.65u l=0.1u
mp4 n3 B1 Y VDD pmos1v w=0.65u l=0.1u
.ends AOI32X1

* Spice subcircuit definition for AOI32X2




.subckt AOI32X2 Y / A0 A1 A2 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 n1 VSS nmos1v w=0.86u l=0.1u
mn2 n1 A2 Y VSS nmos1v w=0.86u l=0.1u
mn3 n2 B0 VSS VSS nmos1v w=0.86u l=0.1u
mn4 n2 B1 Y VSS nmos1v w=0.86u l=0.1u
mp0 n3 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n3 A1 VDD VDD pmos1v w=1.3u l=0.1u
mp2 n3 A2 VDD VDD pmos1v w=1.3u l=0.1u
mp3 n3 B0 Y VDD pmos1v w=1.3u l=0.1u
mp4 n3 B1 Y VDD pmos1v w=1.3u l=0.1u
.ends AOI32X2

* Spice subcircuit definition for AOI32X4




.subckt AOI32X4 Y / A0 A1 A2 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 n1 VSS nmos1v w=1.72u l=0.1u
mn2 n1 A2 Y VSS nmos1v w=1.72u l=0.1u
mn3 n2 B0 VSS VSS nmos1v w=1.72u l=0.1u
mn4 n2 B1 Y VSS nmos1v w=1.72u l=0.1u
mp0 n3 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n3 A1 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n3 A2 VDD VDD pmos1v w=2.6u l=0.1u
mp3 n3 B0 Y VDD pmos1v w=2.6u l=0.1u
mp4 n3 B1 Y VDD pmos1v w=2.6u l=0.1u
.ends AOI32X4

* Spice subcircuit definition for AOI32XL




.subckt AOI32XL Y / A0 A1 A2 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 n1 VSS nmos1v w=0.24u l=0.1u
mn2 n1 A2 Y VSS nmos1v w=0.24u l=0.1u
mn3 n2 B0 VSS VSS nmos1v w=0.24u l=0.1u
mn4 n2 B1 Y VSS nmos1v w=0.24u l=0.1u
mp0 n3 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n3 A1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 A2 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 B0 Y VDD pmos1v w=0.36u l=0.1u
mp4 n3 B1 Y VDD pmos1v w=0.36u l=0.1u
.ends AOI32XL

* Spice subcircuit definition for AOI33X1




.subckt AOI33X1 Y / A0 A1 A2 B0 B1 B2
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 n1 VSS nmos1v w=0.43u l=0.1u
mn2 n1 A2 Y VSS nmos1v w=0.43u l=0.1u
mn3 n2 B0 VSS VSS nmos1v w=0.43u l=0.1u
mn4 n2 B1 n3 VSS nmos1v w=0.43u l=0.1u
mn5 n3 B2 Y VSS nmos1v w=0.43u l=0.1u
mp0 n4 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n4 A1 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n4 A2 VDD VDD pmos1v w=0.65u l=0.1u
mp3 n4 B0 Y VDD pmos1v w=0.65u l=0.1u
mp4 n4 B1 Y VDD pmos1v w=0.65u l=0.1u
mp5 n4 B2 Y VDD pmos1v w=0.65u l=0.1u
.ends AOI33X1

* Spice subcircuit definition for AOI33X2




.subckt AOI33X2 Y / A0 A1 A2 B0 B1 B2
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 n1 VSS nmos1v w=0.86u l=0.1u
mn2 n1 A2 Y VSS nmos1v w=0.86u l=0.1u
mn3 n2 B0 VSS VSS nmos1v w=0.86u l=0.1u
mn4 n2 B1 n3 VSS nmos1v w=0.86u l=0.1u
mn5 n3 B2 Y VSS nmos1v w=0.86u l=0.1u
mp0 n4 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n4 A1 VDD VDD pmos1v w=1.3u l=0.1u
mp2 n4 A2 VDD VDD pmos1v w=1.3u l=0.1u
mp3 n4 B0 Y VDD pmos1v w=1.3u l=0.1u
mp4 n4 B1 Y VDD pmos1v w=1.3u l=0.1u
mp5 n4 B2 Y VDD pmos1v w=1.3u l=0.1u
.ends AOI33X2

* Spice subcircuit definition for AOI33X4




.subckt AOI33X4 Y / A0 A1 A2 B0 B1 B2
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 n1 VSS nmos1v w=1.72u l=0.1u
mn2 n1 A2 Y VSS nmos1v w=1.72u l=0.1u
mn3 n2 B0 VSS VSS nmos1v w=1.72u l=0.1u
mn4 n2 B1 n3 VSS nmos1v w=1.72u l=0.1u
mn5 n3 B2 Y VSS nmos1v w=1.72u l=0.1u
mp0 n4 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n4 A1 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n4 A2 VDD VDD pmos1v w=2.6u l=0.1u
mp3 n4 B0 Y VDD pmos1v w=2.6u l=0.1u
mp4 n4 B1 Y VDD pmos1v w=2.6u l=0.1u
mp5 n4 B2 Y VDD pmos1v w=2.6u l=0.1u
.ends AOI33X4

* Spice subcircuit definition for AOI33XL




.subckt AOI33XL Y / A0 A1 A2 B0 B1 B2
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 n1 VSS nmos1v w=0.24u l=0.1u
mn2 n1 A2 Y VSS nmos1v w=0.24u l=0.1u
mn3 n2 B0 VSS VSS nmos1v w=0.24u l=0.1u
mn4 n2 B1 n3 VSS nmos1v w=0.24u l=0.1u
mn5 n3 B2 Y VSS nmos1v w=0.24u l=0.1u
mp0 n4 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 A2 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 B0 Y VDD pmos1v w=0.36u l=0.1u
mp4 n4 B1 Y VDD pmos1v w=0.36u l=0.1u
mp5 n4 B2 Y VDD pmos1v w=0.36u l=0.1u
.ends AOI33XL

* Spice subcircuit definition for BMXIX2




.subckt BMXIX2 PPN / A M0 M1 S X2
mn0 M0b M0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 M1b M1 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n9 M1 n1 VSS nmos1v w=0.24u l=0.1u
mn11 n0 X2 n2 VSS nmos1v w=0.24u l=0.1u
mn12 n1 X2b n2 VSS nmos1v w=0.24u l=0.1u
mn13 PPN n2 VSS VSS nmos1v w=0.86u l=0.1u
mn2 X2b X2 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 S VSS VSS nmos1v w=0.24u l=0.1u
mn4 n3 M0b n0 VSS nmos1v w=0.24u l=0.1u
mn5 n5 A VSS VSS nmos1v w=0.24u l=0.1u
mn6 n5 M0 n0 VSS nmos1v w=0.24u l=0.1u
mn7 n7 S VSS VSS nmos1v w=0.24u l=0.1u
mn8 n7 M1b n1 VSS nmos1v w=0.24u l=0.1u
mn9 n9 A VSS VSS nmos1v w=0.24u l=0.1u
mp0 M0b M0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 M1b M1 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n10 M1b n1 VDD pmos1v w=0.36u l=0.1u
mp11 n0 X2b n2 VDD pmos1v w=0.36u l=0.1u
mp12 n1 X2 n2 VDD pmos1v w=0.36u l=0.1u
mp13 PPN n2 VDD VDD pmos1v w=1.3u l=0.1u
mp2 X2b X2 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 S VDD VDD pmos1v w=0.36u l=0.1u
mp4 n4 M0 n0 VDD pmos1v w=0.36u l=0.1u
mp5 n6 A VDD VDD pmos1v w=0.36u l=0.1u
mp6 n6 M0b n0 VDD pmos1v w=0.36u l=0.1u
mp7 n8 S VDD VDD pmos1v w=0.36u l=0.1u
mp8 n8 M1 n1 VDD pmos1v w=0.36u l=0.1u
mp9 n10 A VDD VDD pmos1v w=0.36u l=0.1u
.ends BMXIX2

* Spice subcircuit definition for BMXIX4




.subckt BMXIX4 PPN / A M0 M1 S X2
mn0 M0b M0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 M1b M1 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n9 M1 n1 VSS nmos1v w=0.24u l=0.1u
mn11 n0 X2 n2 VSS nmos1v w=0.43u l=0.1u
mn12 n1 X2b n2 VSS nmos1v w=0.43u l=0.1u
mn13 PPN n2 VSS VSS nmos1v w=1.72u l=0.1u
mn2 X2b X2 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 S VSS VSS nmos1v w=0.24u l=0.1u
mn4 n3 M0b n0 VSS nmos1v w=0.24u l=0.1u
mn5 n5 A VSS VSS nmos1v w=0.24u l=0.1u
mn6 n5 M0 n0 VSS nmos1v w=0.24u l=0.1u
mn7 n7 S VSS VSS nmos1v w=0.24u l=0.1u
mn8 n7 M1b n1 VSS nmos1v w=0.24u l=0.1u
mn9 n9 A VSS VSS nmos1v w=0.24u l=0.1u
mp0 M0b M0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 M1b M1 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n10 M1b n1 VDD pmos1v w=0.36u l=0.1u
mp11 n0 X2b n2 VDD pmos1v w=0.65u l=0.1u
mp12 n1 X2 n2 VDD pmos1v w=0.65u l=0.1u
mp13 PPN n2 VDD VDD pmos1v w=2.6u l=0.1u
mp2 X2b X2 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 S VDD VDD pmos1v w=0.36u l=0.1u
mp4 n4 M0 n0 VDD pmos1v w=0.36u l=0.1u
mp5 n6 A VDD VDD pmos1v w=0.36u l=0.1u
mp6 n6 M0b n0 VDD pmos1v w=0.36u l=0.1u
mp7 n8 S VDD VDD pmos1v w=0.36u l=0.1u
mp8 n8 M1 n1 VDD pmos1v w=0.36u l=0.1u
mp9 n10 A VDD VDD pmos1v w=0.36u l=0.1u
.ends BMXIX4

* Spice subcircuit definition for BUFX12




.subckt BUFX12 Y / A
mn0 n0 A VSS VSS nmos1v w=1.29u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=5.16u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.95u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=7.8u l=0.1u
.ends BUFX12

* Spice subcircuit definition for BUFX16




.subckt BUFX16 Y / A
mn0 n0 A VSS VSS nmos1v w=1.72u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=6.88u l=0.1u
mp0 n0 A VDD VDD pmos1v w=2.6u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=10.4u l=0.1u
.ends BUFX16

* Spice subcircuit definition for BUFX2




.subckt BUFX2 Y / A
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends BUFX2

* Spice subcircuit definition for BUFX20




.subckt BUFX20 Y / A
mn0 n0 A VSS VSS nmos1v w=2.15u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=8.6u l=0.1u
mp0 n0 A VDD VDD pmos1v w=3.25u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=13.0u l=0.1u
.ends BUFX20

* Spice subcircuit definition for BUFX3




.subckt BUFX3 Y / A
mn0 n0 A VSS VSS nmos1v w=0.43u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=1.29u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=1.95u l=0.1u
.ends BUFX3

* Spice subcircuit definition for BUFX4




.subckt BUFX4 Y / A
mn0 n0 A VSS VSS nmos1v w=0.43u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends BUFX4

* Spice subcircuit definition for BUFX6




.subckt BUFX6 Y / A
mn0 n0 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=2.58u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=3.9u l=0.1u
.ends BUFX6

* Spice subcircuit definition for BUFX8




.subckt BUFX8 Y / A
mn0 n0 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=3.44u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=5.2u l=0.1u
.ends BUFX8

* Spice subcircuit definition for CLKAND2X12




.subckt CLKAND2X12 Y / A B
mn0 n1 A VSS VSS nmos1v w=2.58u l=0.1u
mn1 n1 B n0 VSS nmos1v w=2.58u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=5.16u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.95u l=0.1u
mp1 n0 B VDD VDD pmos1v w=1.95u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=7.8u l=0.1u
.ends CLKAND2X12

* Spice subcircuit definition for CLKAND2X2




.subckt CLKAND2X2 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.48u l=0.1u
mn1 n1 B n0 VSS nmos1v w=0.48u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends CLKAND2X2

* Spice subcircuit definition for CLKAND2X3




.subckt CLKAND2X3 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n1 B n0 VSS nmos1v w=0.86u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=1.29u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 n0 B VDD VDD pmos1v w=0.65u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=1.95u l=0.1u
.ends CLKAND2X3

* Spice subcircuit definition for CLKAND2X4




.subckt CLKAND2X4 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n1 B n0 VSS nmos1v w=0.86u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 n0 B VDD VDD pmos1v w=0.65u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends CLKAND2X4

* Spice subcircuit definition for CLKAND2X6




.subckt CLKAND2X6 Y / A B
mn0 n1 A VSS VSS nmos1v w=1.72u l=0.1u
mn1 n1 B n0 VSS nmos1v w=1.72u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=2.58u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n0 B VDD VDD pmos1v w=1.3u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=3.9u l=0.1u
.ends CLKAND2X6

* Spice subcircuit definition for CLKAND2X8




.subckt CLKAND2X8 Y / A B
mn0 n1 A VSS VSS nmos1v w=1.72u l=0.1u
mn1 n1 B n0 VSS nmos1v w=1.72u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=3.44u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n0 B VDD VDD pmos1v w=1.3u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=5.2u l=0.1u
.ends CLKAND2X8

* Spice subcircuit definition for CLKBUFX12




.subckt CLKBUFX12 Y / A
mn0 n0 A VSS VSS nmos1v w=1.29u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=5.16u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.95u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=7.8u l=0.1u
.ends CLKBUFX12

* Spice subcircuit definition for CLKBUFX16




.subckt CLKBUFX16 Y / A
mn0 n0 A VSS VSS nmos1v w=1.72u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=6.88u l=0.1u
mp0 n0 A VDD VDD pmos1v w=2.6u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=10.4u l=0.1u
.ends CLKBUFX16

* Spice subcircuit definition for CLKBUFX2




.subckt CLKBUFX2 Y / A
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends CLKBUFX2

* Spice subcircuit definition for CLKBUFX20




.subckt CLKBUFX20 Y / A
mn0 n0 A VSS VSS nmos1v w=2.15u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=8.6u l=0.1u
mp0 n0 A VDD VDD pmos1v w=3.25u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=13.0u l=0.1u
.ends CLKBUFX20

* Spice subcircuit definition for CLKBUFX3




.subckt CLKBUFX3 Y / A
mn0 n0 A VSS VSS nmos1v w=0.43u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=1.29u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=1.95u l=0.1u
.ends CLKBUFX3

* Spice subcircuit definition for CLKBUFX4




.subckt CLKBUFX4 Y / A
mn0 n0 A VSS VSS nmos1v w=0.43u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends CLKBUFX4

* Spice subcircuit definition for CLKBUFX6




.subckt CLKBUFX6 Y / A
mn0 n0 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=2.58u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=3.9u l=0.1u
.ends CLKBUFX6

* Spice subcircuit definition for CLKBUFX8




.subckt CLKBUFX8 Y / A
mn0 n0 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=3.44u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=5.2u l=0.1u
.ends CLKBUFX8

* Spice subcircuit definition for CLKINVX1




.subckt CLKINVX1 Y / A
mn0 Y A VSS VSS nmos1v w=0.43u l=0.1u
mp0 Y A VDD VDD pmos1v w=0.65u l=0.1u
.ends CLKINVX1

* Spice subcircuit definition for CLKINVX12




.subckt CLKINVX12 Y / A
mn0 Y A VSS VSS nmos1v w=5.16u l=0.1u
mp0 Y A VDD VDD pmos1v w=7.8u l=0.1u
.ends CLKINVX12

* Spice subcircuit definition for CLKINVX16




.subckt CLKINVX16 Y / A
mn0 Y A VSS VSS nmos1v w=6.88u l=0.1u
mp0 Y A VDD VDD pmos1v w=10.4u l=0.1u
.ends CLKINVX16

* Spice subcircuit definition for CLKINVX2




.subckt CLKINVX2 Y / A
mn0 Y A VSS VSS nmos1v w=0.86u l=0.1u
mp0 Y A VDD VDD pmos1v w=1.3u l=0.1u
.ends CLKINVX2

* Spice subcircuit definition for CLKINVX20




.subckt CLKINVX20 Y / A
mn0 Y A VSS VSS nmos1v w=8.6u l=0.1u
mp0 Y A VDD VDD pmos1v w=13.0u l=0.1u
.ends CLKINVX20

* Spice subcircuit definition for CLKINVX3




.subckt CLKINVX3 Y / A
mn0 Y A VSS VSS nmos1v w=1.29u l=0.1u
mp0 Y A VDD VDD pmos1v w=1.95u l=0.1u
.ends CLKINVX3

* Spice subcircuit definition for CLKINVX4




.subckt CLKINVX4 Y / A
mn0 Y A VSS VSS nmos1v w=1.72u l=0.1u
mp0 Y A VDD VDD pmos1v w=2.6u l=0.1u
.ends CLKINVX4

* Spice subcircuit definition for CLKINVX6




.subckt CLKINVX6 Y / A
mn0 Y A VSS VSS nmos1v w=2.58u l=0.1u
mp0 Y A VDD VDD pmos1v w=3.9u l=0.1u
.ends CLKINVX6

* Spice subcircuit definition for CLKINVX8




.subckt CLKINVX8 Y / A
mn0 Y A VSS VSS nmos1v w=3.44u l=0.1u
mp0 Y A VDD VDD pmos1v w=5.2u l=0.1u
.ends CLKINVX8

* Spice subcircuit definition for CLKMX2X12




.subckt CLKMX2X12 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.34u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.34u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.34u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.34u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=5.16u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.52u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.52u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.52u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.52u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=7.8u l=0.1u
.ends CLKMX2X12

* Spice subcircuit definition for CLKMX2X2




.subckt CLKMX2X2 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends CLKMX2X2

* Spice subcircuit definition for CLKMX2X3




.subckt CLKMX2X3 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.43u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.43u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.43u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.43u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=1.29u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.65u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.65u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.65u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.65u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=1.95u l=0.1u
.ends CLKMX2X3

* Spice subcircuit definition for CLKMX2X4




.subckt CLKMX2X4 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.34u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.34u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.34u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.34u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.52u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.52u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.52u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.52u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends CLKMX2X4

* Spice subcircuit definition for CLKMX2X6




.subckt CLKMX2X6 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.34u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.34u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.34u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.34u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=2.58u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.52u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.52u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.52u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.52u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=3.9u l=0.1u
.ends CLKMX2X6

* Spice subcircuit definition for CLKMX2X8




.subckt CLKMX2X8 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.34u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.34u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.34u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.34u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=3.44u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.52u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.52u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.52u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.52u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=5.2u l=0.1u
.ends CLKMX2X8

* Spice subcircuit definition for CLKXOR2X1




.subckt CLKXOR2X1 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n2 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 B n0 VSS nmos1v w=0.24u l=0.1u
mn4 n1 n2 n0 VSS nmos1v w=0.24u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 n2 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n1 B n0 VDD pmos1v w=0.36u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends CLKXOR2X1

* Spice subcircuit definition for CLKXOR2X2




.subckt CLKXOR2X2 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n2 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 B n0 VSS nmos1v w=0.24u l=0.1u
mn4 n1 n2 n0 VSS nmos1v w=0.24u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 n2 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n1 B n0 VDD pmos1v w=0.36u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends CLKXOR2X2

* Spice subcircuit definition for CLKXOR2X4




.subckt CLKXOR2X4 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n2 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 n1 VSS VSS nmos1v w=0.34u l=0.1u
mn3 n3 B n0 VSS nmos1v w=0.34u l=0.1u
mn4 n1 n2 n0 VSS nmos1v w=0.34u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 n1 VDD VDD pmos1v w=0.52u l=0.1u
mp3 n4 n2 n0 VDD pmos1v w=0.52u l=0.1u
mp4 n1 B n0 VDD pmos1v w=0.52u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends CLKXOR2X4

* Spice subcircuit definition for CLKXOR2X8




.subckt CLKXOR2X8 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n2 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 n1 VSS VSS nmos1v w=0.34u l=0.1u
mn3 n3 B n0 VSS nmos1v w=0.34u l=0.1u
mn4 n1 n2 n0 VSS nmos1v w=0.34u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=3.44u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 n1 VDD VDD pmos1v w=0.52u l=0.1u
mp3 n4 n2 n0 VDD pmos1v w=0.52u l=0.1u
mp4 n1 B n0 VDD pmos1v w=0.52u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=5.2u l=0.1u
.ends CLKXOR2X8

* Spice subcircuit definition for DFFHQX1




.subckt DFFHQX1 Q / CK D
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
.ends DFFHQX1

* Spice subcircuit definition for DFFHQX2




.subckt DFFHQX2 Q / CK D
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
.ends DFFHQX2

* Spice subcircuit definition for DFFHQX4




.subckt DFFHQX4 Q / CK D
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
.ends DFFHQX4

* Spice subcircuit definition for DFFHQX8




.subckt DFFHQX8 Q / CK D
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=1.29u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=3.44u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.95u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=5.2u l=0.1u
.ends DFFHQX8

* Spice subcircuit definition for DFFNSRX1




.subckt DFFNSRX1 Q QN / CKN D RN SN
mn20 CKNb CKN VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKNbb CKNb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKNbb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKNb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKNb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKNbb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mp20 CKNb CKN VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKNbb CKNb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKNb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKNbb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKNbb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKNb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
.ends DFFNSRX1

* Spice subcircuit definition for DFFNSRX2




.subckt DFFNSRX2 Q QN / CKN D RN SN
mn20 CKNb CKN VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKNbb CKNb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKNbb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKNb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKNb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKNbb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mp20 CKNb CKN VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKNbb CKNb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKNb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKNbb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKNbb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKNb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
.ends DFFNSRX2

* Spice subcircuit definition for DFFNSRX4




.subckt DFFNSRX4 Q QN / CKN D RN SN
mn20 CKNb CKN VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKNbb CKNb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKNbb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKNb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKNb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKNbb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mp20 CKNb CKN VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKNbb CKNb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKNb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKNbb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKNbb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKNb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
.ends DFFNSRX4

* Spice subcircuit definition for DFFNSRXL




.subckt DFFNSRXL Q QN / CKN D RN SN
mn20 CKNb CKN VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKNbb CKNb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKNbb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKNb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKNb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKNbb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mp20 CKNb CKN VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKNbb CKNb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKNb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKNbb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKNbb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKNb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
.ends DFFNSRXL

* Spice subcircuit definition for DFFQX1




.subckt DFFQX1 Q / CK D
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
.ends DFFQX1

* Spice subcircuit definition for DFFQX2




.subckt DFFQX2 Q / CK D
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
.ends DFFQX2

* Spice subcircuit definition for DFFQX4




.subckt DFFQX4 Q / CK D
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
.ends DFFQX4

* Spice subcircuit definition for DFFQXL




.subckt DFFQXL Q / CK D
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
.ends DFFQXL

* Spice subcircuit definition for DFFRHQX1




.subckt DFFRHQX1 Q / CK D RN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.34u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.34u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=0.34u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=0.34u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=0.52u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
.ends DFFRHQX1

* Spice subcircuit definition for DFFRHQX2




.subckt DFFRHQX2 Q / CK D RN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.34u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.34u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=0.34u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=0.34u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=0.52u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
.ends DFFRHQX2

* Spice subcircuit definition for DFFRHQX4




.subckt DFFRHQX4 Q / CK D RN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.34u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.34u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=0.68u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=0.68u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=1.04u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
.ends DFFRHQX4

* Spice subcircuit definition for DFFRHQX8




.subckt DFFRHQX8 Q / CK D RN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.34u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.34u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=1.29u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=1.29u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=3.44u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=1.95u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=1.95u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=5.2u l=0.1u
.ends DFFRHQX8

* Spice subcircuit definition for DFFRX1




.subckt DFFRX1 Q QN / CK D RN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.24u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.24u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=0.24u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=0.24u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=0.36u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
.ends DFFRX1

* Spice subcircuit definition for DFFRX2




.subckt DFFRX2 Q QN / CK D RN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.24u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.24u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=0.34u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=0.34u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=0.52u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
.ends DFFRX2

* Spice subcircuit definition for DFFRX4




.subckt DFFRX4 Q QN / CK D RN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.24u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.24u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=0.68u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=0.68u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=1.04u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
.ends DFFRX4

* Spice subcircuit definition for DFFRXL




.subckt DFFRXL Q QN / CK D RN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.24u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.24u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=0.24u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=0.24u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=0.36u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
.ends DFFRXL

* Spice subcircuit definition for DFFSHQX1




.subckt DFFSHQX1 Q / CK D SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
.ends DFFSHQX1

* Spice subcircuit definition for DFFSHQX2




.subckt DFFSHQX2 Q / CK D SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
.ends DFFSHQX2

* Spice subcircuit definition for DFFSHQX4




.subckt DFFSHQX4 Q / CK D SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
.ends DFFSHQX4

* Spice subcircuit definition for DFFSHQX8




.subckt DFFSHQX8 Q / CK D SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=1.29u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=3.44u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=1.95u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=5.2u l=0.1u
.ends DFFSHQX8

* Spice subcircuit definition for DFFSRHQX1




.subckt DFFSRHQX1 Q / CK D RN SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.34u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.34u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.52u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
.ends DFFSRHQX1

* Spice subcircuit definition for DFFSRHQX2




.subckt DFFSRHQX2 Q / CK D RN SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.34u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.34u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.52u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
.ends DFFSRHQX2

* Spice subcircuit definition for DFFSRHQX4




.subckt DFFSRHQX4 Q / CK D RN SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.34u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.34u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.52u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
.ends DFFSRHQX4

* Spice subcircuit definition for DFFSRHQX8




.subckt DFFSRHQX8 Q / CK D RN SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.34u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.34u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=1.29u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.34u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=3.44u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.52u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=1.95u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.52u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=5.2u l=0.1u
.ends DFFSRHQX8

* Spice subcircuit definition for DFFSRX1




.subckt DFFSRX1 Q QN / CK D RN SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
.ends DFFSRX1

* Spice subcircuit definition for DFFSRX2




.subckt DFFSRX2 Q QN / CK D RN SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
.ends DFFSRX2

* Spice subcircuit definition for DFFSRX4




.subckt DFFSRX4 Q QN / CK D RN SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
.ends DFFSRX4

* Spice subcircuit definition for DFFSRXL




.subckt DFFSRXL Q QN / CK D RN SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
.ends DFFSRXL

* Spice subcircuit definition for DFFSX1




.subckt DFFSX1 Q QN / CK D SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
.ends DFFSX1

* Spice subcircuit definition for DFFSX2




.subckt DFFSX2 Q QN / CK D SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
.ends DFFSX2

* Spice subcircuit definition for DFFSX4




.subckt DFFSX4 Q QN / CK D SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
.ends DFFSX4

* Spice subcircuit definition for DFFSXL




.subckt DFFSXL Q QN / CK D SN
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
.ends DFFSXL

* Spice subcircuit definition for DFFTRX1




.subckt DFFTRX1 Q QN / CK D RN
mn0 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 D Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mp0 Db RN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
.ends DFFTRX1

* Spice subcircuit definition for DFFTRX2




.subckt DFFTRX2 Q QN / CK D RN
mn0 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 D Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mp0 Db RN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
.ends DFFTRX2

* Spice subcircuit definition for DFFTRX4




.subckt DFFTRX4 Q QN / CK D RN
mn0 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 D Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mp0 Db RN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
.ends DFFTRX4

* Spice subcircuit definition for DFFTRXL




.subckt DFFTRXL Q QN / CK D RN
mn0 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 D Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mp0 Db RN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
.ends DFFTRXL

* Spice subcircuit definition for DFFX1




.subckt DFFX1 Q QN / CK D
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
.ends DFFX1

* Spice subcircuit definition for DFFX2




.subckt DFFX2 Q QN / CK D
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
.ends DFFX2

* Spice subcircuit definition for DFFX4




.subckt DFFX4 Q QN / CK D
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
.ends DFFX4

* Spice subcircuit definition for DFFXL




.subckt DFFXL Q QN / CK D
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 D VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 D VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
.ends DFFXL

* Spice subcircuit definition for DLY1X1




.subckt DLY1X1 Y / A
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n4 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n4 VDD n1 VSS nmos1v w=0.24u l=0.1u
mn3 n2 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn4 Y n2 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n5 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n5 VSS n1 VDD pmos1v w=0.36u l=0.1u
mp3 n2 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp4 Y n2 VDD VDD pmos1v w=0.65u l=0.1u
.ends DLY1X1

* Spice subcircuit definition for DLY1X4




.subckt DLY1X4 Y / A
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n4 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n4 VDD n1 VSS nmos1v w=0.24u l=0.1u
mn3 n2 n1 VSS VSS nmos1v w=0.43u l=0.1u
mn4 Y n2 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n5 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n5 VSS n1 VDD pmos1v w=0.36u l=0.1u
mp3 n2 n1 VDD VDD pmos1v w=0.65u l=0.1u
mp4 Y n2 VDD VDD pmos1v w=2.6u l=0.1u
.ends DLY1X4

* Spice subcircuit definition for DLY2X1




.subckt DLY2X1 Y / A
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n6 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n6 VDD n1 VSS nmos1v w=0.24u l=0.1u
mn3 n8 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn4 n8 VDD n2 VSS nmos1v w=0.24u l=0.1u
mn5 n10 n2 VSS VSS nmos1v w=0.24u l=0.1u
mn6 n10 VDD n3 VSS nmos1v w=0.24u l=0.1u
mn7 n4 n3 VSS VSS nmos1v w=0.24u l=0.1u
mn8 Y n4 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n7 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n7 VSS n1 VDD pmos1v w=0.36u l=0.1u
mp3 n9 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp4 n9 VSS n2 VDD pmos1v w=0.36u l=0.1u
mp5 n11 n2 VDD VDD pmos1v w=0.36u l=0.1u
mp6 n11 VSS n3 VDD pmos1v w=0.36u l=0.1u
mp7 n4 n3 VDD VDD pmos1v w=0.36u l=0.1u
mp8 Y n4 VDD VDD pmos1v w=0.65u l=0.1u
.ends DLY2X1

* Spice subcircuit definition for DLY2X4




.subckt DLY2X4 Y / A
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n6 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n6 VDD n1 VSS nmos1v w=0.24u l=0.1u
mn3 n8 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn4 n8 VDD n2 VSS nmos1v w=0.24u l=0.1u
mn5 n10 n2 VSS VSS nmos1v w=0.24u l=0.1u
mn6 n10 VDD n3 VSS nmos1v w=0.24u l=0.1u
mn7 n4 n3 VSS VSS nmos1v w=0.43u l=0.1u
mn8 Y n4 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n7 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n7 VSS n1 VDD pmos1v w=0.36u l=0.1u
mp3 n9 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp4 n9 VSS n2 VDD pmos1v w=0.36u l=0.1u
mp5 n11 n2 VDD VDD pmos1v w=0.36u l=0.1u
mp6 n11 VSS n3 VDD pmos1v w=0.36u l=0.1u
mp7 n4 n3 VDD VDD pmos1v w=0.65u l=0.1u
mp8 Y n4 VDD VDD pmos1v w=2.6u l=0.1u
.ends DLY2X4

* Spice subcircuit definition for DLY3X1




.subckt DLY3X1 Y / A
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n8 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n16 VDD n5 VSS nmos1v w=0.24u l=0.1u
mn11 n6 n5 VSS VSS nmos1v w=0.24u l=0.1u
mn12 Y n6 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n8 VDD n1 VSS nmos1v w=0.24u l=0.1u
mn3 n10 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn4 n10 VDD n2 VSS nmos1v w=0.24u l=0.1u
mn5 n12 n2 VSS VSS nmos1v w=0.24u l=0.1u
mn6 n12 VDD n3 VSS nmos1v w=0.24u l=0.1u
mn7 n14 n3 VSS VSS nmos1v w=0.24u l=0.1u
mn8 n14 VDD n4 VSS nmos1v w=0.24u l=0.1u
mn9 n16 n4 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n9 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n17 VSS n5 VDD pmos1v w=0.36u l=0.1u
mp11 n6 n5 VDD VDD pmos1v w=0.36u l=0.1u
mp12 Y n6 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n9 VSS n1 VDD pmos1v w=0.36u l=0.1u
mp3 n11 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp4 n11 VSS n2 VDD pmos1v w=0.36u l=0.1u
mp5 n13 n2 VDD VDD pmos1v w=0.36u l=0.1u
mp6 n13 VSS n3 VDD pmos1v w=0.36u l=0.1u
mp7 n15 n3 VDD VDD pmos1v w=0.36u l=0.1u
mp8 n15 VSS n4 VDD pmos1v w=0.36u l=0.1u
mp9 n17 n4 VDD VDD pmos1v w=0.36u l=0.1u
.ends DLY3X1

* Spice subcircuit definition for DLY3X4




.subckt DLY3X4 Y / A
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n8 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n16 VDD n5 VSS nmos1v w=0.24u l=0.1u
mn11 n6 n5 VSS VSS nmos1v w=0.43u l=0.1u
mn12 Y n6 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n8 VDD n1 VSS nmos1v w=0.24u l=0.1u
mn3 n10 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn4 n10 VDD n2 VSS nmos1v w=0.24u l=0.1u
mn5 n12 n2 VSS VSS nmos1v w=0.24u l=0.1u
mn6 n12 VDD n3 VSS nmos1v w=0.24u l=0.1u
mn7 n14 n3 VSS VSS nmos1v w=0.24u l=0.1u
mn8 n14 VDD n4 VSS nmos1v w=0.24u l=0.1u
mn9 n16 n4 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n9 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n17 VSS n5 VDD pmos1v w=0.36u l=0.1u
mp11 n6 n5 VDD VDD pmos1v w=0.65u l=0.1u
mp12 Y n6 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n9 VSS n1 VDD pmos1v w=0.36u l=0.1u
mp3 n11 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp4 n11 VSS n2 VDD pmos1v w=0.36u l=0.1u
mp5 n13 n2 VDD VDD pmos1v w=0.36u l=0.1u
mp6 n13 VSS n3 VDD pmos1v w=0.36u l=0.1u
mp7 n15 n3 VDD VDD pmos1v w=0.36u l=0.1u
mp8 n15 VSS n4 VDD pmos1v w=0.36u l=0.1u
mp9 n17 n4 VDD VDD pmos1v w=0.36u l=0.1u
.ends DLY3X4

* Spice subcircuit definition for DLY4X1




.subckt DLY4X1 Y / A
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n10 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n18 VDD n5 VSS nmos1v w=0.24u l=0.1u
mn11 n20 n5 VSS VSS nmos1v w=0.24u l=0.1u
mn12 n20 VDD n6 VSS nmos1v w=0.24u l=0.1u
mn13 n22 n6 VSS VSS nmos1v w=0.24u l=0.1u
mn14 n22 VDD n7 VSS nmos1v w=0.24u l=0.1u
mn15 n8 n7 VSS VSS nmos1v w=0.24u l=0.1u
mn16 Y n8 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n10 VDD n1 VSS nmos1v w=0.24u l=0.1u
mn3 n12 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn4 n12 VDD n2 VSS nmos1v w=0.24u l=0.1u
mn5 n14 n2 VSS VSS nmos1v w=0.24u l=0.1u
mn6 n14 VDD n3 VSS nmos1v w=0.24u l=0.1u
mn7 n16 n3 VSS VSS nmos1v w=0.24u l=0.1u
mn8 n16 VDD n4 VSS nmos1v w=0.24u l=0.1u
mn9 n18 n4 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n11 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n19 VSS n5 VDD pmos1v w=0.36u l=0.1u
mp11 n21 n5 VDD VDD pmos1v w=0.36u l=0.1u
mp12 n21 VSS n6 VDD pmos1v w=0.36u l=0.1u
mp13 n23 n6 VDD VDD pmos1v w=0.36u l=0.1u
mp14 n23 VSS n7 VDD pmos1v w=0.36u l=0.1u
mp15 n8 n7 VDD VDD pmos1v w=0.36u l=0.1u
mp16 Y n8 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n11 VSS n1 VDD pmos1v w=0.36u l=0.1u
mp3 n13 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp4 n13 VSS n2 VDD pmos1v w=0.36u l=0.1u
mp5 n15 n2 VDD VDD pmos1v w=0.36u l=0.1u
mp6 n15 VSS n3 VDD pmos1v w=0.36u l=0.1u
mp7 n17 n3 VDD VDD pmos1v w=0.36u l=0.1u
mp8 n17 VSS n4 VDD pmos1v w=0.36u l=0.1u
mp9 n19 n4 VDD VDD pmos1v w=0.36u l=0.1u
.ends DLY4X1

* Spice subcircuit definition for DLY4X4




.subckt DLY4X4 Y / A
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n10 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n18 VDD n5 VSS nmos1v w=0.24u l=0.1u
mn11 n20 n5 VSS VSS nmos1v w=0.24u l=0.1u
mn12 n20 VDD n6 VSS nmos1v w=0.24u l=0.1u
mn13 n22 n6 VSS VSS nmos1v w=0.24u l=0.1u
mn14 n22 VDD n7 VSS nmos1v w=0.24u l=0.1u
mn15 n8 n7 VSS VSS nmos1v w=0.43u l=0.1u
mn16 Y n8 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n10 VDD n1 VSS nmos1v w=0.24u l=0.1u
mn3 n12 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn4 n12 VDD n2 VSS nmos1v w=0.24u l=0.1u
mn5 n14 n2 VSS VSS nmos1v w=0.24u l=0.1u
mn6 n14 VDD n3 VSS nmos1v w=0.24u l=0.1u
mn7 n16 n3 VSS VSS nmos1v w=0.24u l=0.1u
mn8 n16 VDD n4 VSS nmos1v w=0.24u l=0.1u
mn9 n18 n4 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n11 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n19 VSS n5 VDD pmos1v w=0.36u l=0.1u
mp11 n21 n5 VDD VDD pmos1v w=0.36u l=0.1u
mp12 n21 VSS n6 VDD pmos1v w=0.36u l=0.1u
mp13 n23 n6 VDD VDD pmos1v w=0.36u l=0.1u
mp14 n23 VSS n7 VDD pmos1v w=0.36u l=0.1u
mp15 n8 n7 VDD VDD pmos1v w=0.65u l=0.1u
mp16 Y n8 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n11 VSS n1 VDD pmos1v w=0.36u l=0.1u
mp3 n13 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp4 n13 VSS n2 VDD pmos1v w=0.36u l=0.1u
mp5 n15 n2 VDD VDD pmos1v w=0.36u l=0.1u
mp6 n15 VSS n3 VDD pmos1v w=0.36u l=0.1u
mp7 n17 n3 VDD VDD pmos1v w=0.36u l=0.1u
mp8 n17 VSS n4 VDD pmos1v w=0.36u l=0.1u
mp9 n19 n4 VDD VDD pmos1v w=0.36u l=0.1u
.ends DLY4X4

* Spice subcircuit definition for EDFFHQX1




.subckt EDFFHQX1 Q / CK D E
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 qbint Eb Db VSS nmos1v w=0.43u l=0.1u
mn2 n0 D VSS VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn3 n0 E Db VSS nmos1v w=0.43u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 qbint E Db VDD pmos1v w=0.65u l=0.1u
mp2 n1 D VDD VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp3 n1 Eb Db VDD pmos1v w=0.65u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
.ends EDFFHQX1

* Spice subcircuit definition for EDFFHQX2




.subckt EDFFHQX2 Q / CK D E
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 qbint Eb Db VSS nmos1v w=0.43u l=0.1u
mn2 n0 D VSS VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn3 n0 E Db VSS nmos1v w=0.43u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.43u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 qbint E Db VDD pmos1v w=0.65u l=0.1u
mp2 n1 D VDD VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp3 n1 Eb Db VDD pmos1v w=0.65u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.65u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
.ends EDFFHQX2

* Spice subcircuit definition for EDFFHQX4




.subckt EDFFHQX4 Q / CK D E
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 qbint Eb Db VSS nmos1v w=0.43u l=0.1u
mn2 n0 D VSS VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn3 n0 E Db VSS nmos1v w=0.43u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 qbint E Db VDD pmos1v w=0.65u l=0.1u
mp2 n1 D VDD VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp3 n1 Eb Db VDD pmos1v w=0.65u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
.ends EDFFHQX4

* Spice subcircuit definition for EDFFHQX8




.subckt EDFFHQX8 Q / CK D E
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 qbint Eb Db VSS nmos1v w=0.43u l=0.1u
mn2 n0 D VSS VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn3 n0 E Db VSS nmos1v w=0.43u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=1.29u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=3.44u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 qbint E Db VDD pmos1v w=0.65u l=0.1u
mp2 n1 D VDD VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp3 n1 Eb Db VDD pmos1v w=0.65u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.95u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=5.2u l=0.1u
.ends EDFFHQX8

* Spice subcircuit definition for EDFFTRX1




.subckt EDFFTRX1 Q QN / CK D E RN
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 Db D VSS VSS nmos1v w=0.24u l=0.1u
mn2 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 Dp VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 Dp RNb VSS VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn4 n0 Eb VSS VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn5 n0 qbint Dp VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mn6 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn7 n1 Db Dp VSS nmos1v w=0.24u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp2 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 Dp VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n2 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp4 n2 Eb n3 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp5 n2 qbint n3 VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
mp6 n3 E Dp VDD pmos1v w=0.36u l=0.1u
mp7 n3 Db Dp VDD pmos1v w=0.36u l=0.1u
.ends EDFFTRX1

* Spice subcircuit definition for EDFFTRX2




.subckt EDFFTRX2 Q QN / CK D E RN
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 Db D VSS VSS nmos1v w=0.24u l=0.1u
mn2 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 Dp VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 Dp RNb VSS VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn4 n0 Eb VSS VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.43u l=0.1u
mn5 n0 qbint Dp VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mn6 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn7 n1 Db Dp VSS nmos1v w=0.24u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp2 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 Dp VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n2 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp4 n2 Eb n3 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.65u l=0.1u
mp5 n2 qbint n3 VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
mp6 n3 E Dp VDD pmos1v w=0.36u l=0.1u
mp7 n3 Db Dp VDD pmos1v w=0.36u l=0.1u
.ends EDFFTRX2

* Spice subcircuit definition for EDFFTRX4




.subckt EDFFTRX4 Q QN / CK D E RN
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 Db D VSS VSS nmos1v w=0.24u l=0.1u
mn2 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 Dp VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 Dp RNb VSS VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn4 n0 Eb VSS VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn5 n0 qbint Dp VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mn6 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn7 n1 Db Dp VSS nmos1v w=0.24u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp2 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 Dp VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n2 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp4 n2 Eb n3 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp5 n2 qbint n3 VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
mp6 n3 E Dp VDD pmos1v w=0.36u l=0.1u
mp7 n3 Db Dp VDD pmos1v w=0.36u l=0.1u
.ends EDFFTRX4

* Spice subcircuit definition for EDFFTRXL




.subckt EDFFTRXL Q QN / CK D E RN
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 Db D VSS VSS nmos1v w=0.24u l=0.1u
mn2 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 n21 Dp VSS VSS nmos1v w=0.24u l=0.1u
mn26 n21 CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 Dp RNb VSS VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn4 n0 Eb VSS VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn5 n0 qbint Dp VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn7 n1 Db Dp VSS nmos1v w=0.24u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp2 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 n22 Dp VDD VDD pmos1v w=0.36u l=0.1u
mp26 n22 CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n2 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp4 n2 Eb n3 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp5 n2 qbint n3 VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
mp6 n3 E Dp VDD pmos1v w=0.36u l=0.1u
mp7 n3 Db Dp VDD pmos1v w=0.36u l=0.1u
.ends EDFFTRXL

* Spice subcircuit definition for EDFFX1




.subckt EDFFX1 Q QN / CK D E
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 qbint Eb Db VSS nmos1v w=0.24u l=0.1u
mn2 n0 D VSS VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 n0 E Db VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 qbint E Db VDD pmos1v w=0.36u l=0.1u
mp2 n1 D VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n1 Eb Db VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
.ends EDFFX1

* Spice subcircuit definition for EDFFX2




.subckt EDFFX2 Q QN / CK D E
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 qbint Eb Db VSS nmos1v w=0.24u l=0.1u
mn2 n0 D VSS VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 n0 E Db VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.43u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 qbint E Db VDD pmos1v w=0.36u l=0.1u
mp2 n1 D VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n1 Eb Db VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.65u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
.ends EDFFX2

* Spice subcircuit definition for EDFFX4




.subckt EDFFX4 Q QN / CK D E
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 qbint Eb Db VSS nmos1v w=0.24u l=0.1u
mn2 n0 D VSS VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 n0 E Db VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 qbint E Db VDD pmos1v w=0.36u l=0.1u
mp2 n1 D VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n1 Eb Db VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
.ends EDFFX4

* Spice subcircuit definition for EDFFXL




.subckt EDFFXL Q QN / CK D E
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 qbint Eb Db VSS nmos1v w=0.24u l=0.1u
mn2 n0 D VSS VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 n0 E Db VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 qbint E Db VDD pmos1v w=0.36u l=0.1u
mp2 n1 D VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n1 Eb Db VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
.ends EDFFXL

* Spice subcircuit definition for HOLDX1




.subckt HOLDX1 Y
mn0 n0 Y VSS VSS nmos1v w=0.43u l=0.1u
mn1 nn1 n0 Y VSS nmos1v w=0.24u l=0.1u
mn2 nn2 n0 nn1 VSS nmos1v w=0.24u l=0.1u
mn3 nn2 n0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 Y VDD VDD pmos1v w=0.65u l=0.1u
mp1 np1 n0 Y VDD pmos1v w=0.36u l=0.1u
mp2 np2 n0 np1 VDD pmos1v w=0.36u l=0.1u
mp3 np2 n0 VDD VDD pmos1v w=0.36u l=0.1u
.ends HOLDX1

* Spice subcircuit definition for INVX1




.subckt INVX1 Y / A
mn0 Y A VSS VSS nmos1v w=0.43u l=0.1u
mp0 Y A VDD VDD pmos1v w=0.65u l=0.1u
.ends INVX1

* Spice subcircuit definition for INVX12




.subckt INVX12 Y / A
mn0 Y A VSS VSS nmos1v w=5.16u l=0.1u
mp0 Y A VDD VDD pmos1v w=7.8u l=0.1u
.ends INVX12

* Spice subcircuit definition for INVX16




.subckt INVX16 Y / A
mn0 Y A VSS VSS nmos1v w=6.88u l=0.1u
mp0 Y A VDD VDD pmos1v w=10.4u l=0.1u
.ends INVX16

* Spice subcircuit definition for INVX2




.subckt INVX2 Y / A
mn0 Y A VSS VSS nmos1v w=0.86u l=0.1u
mp0 Y A VDD VDD pmos1v w=1.3u l=0.1u
.ends INVX2

* Spice subcircuit definition for INVX20




.subckt INVX20 Y / A
mn0 Y A VSS VSS nmos1v w=8.6u l=0.1u
mp0 Y A VDD VDD pmos1v w=13.0u l=0.1u
.ends INVX20

* Spice subcircuit definition for INVX3




.subckt INVX3 Y / A
mn0 Y A VSS VSS nmos1v w=1.29u l=0.1u
mp0 Y A VDD VDD pmos1v w=1.95u l=0.1u
.ends INVX3

* Spice subcircuit definition for INVX4




.subckt INVX4 Y / A
mn0 Y A VSS VSS nmos1v w=1.72u l=0.1u
mp0 Y A VDD VDD pmos1v w=2.6u l=0.1u
.ends INVX4

* Spice subcircuit definition for INVX6




.subckt INVX6 Y / A
mn0 Y A VSS VSS nmos1v w=2.58u l=0.1u
mp0 Y A VDD VDD pmos1v w=3.9u l=0.1u
.ends INVX6

* Spice subcircuit definition for INVX8




.subckt INVX8 Y / A
mn0 Y A VSS VSS nmos1v w=3.44u l=0.1u
mp0 Y A VDD VDD pmos1v w=5.2u l=0.1u
.ends INVX8

* Spice subcircuit definition for INVXL




.subckt INVXL Y / A
mn0 Y A VSS VSS nmos1v w=0.24u l=0.1u
mp0 Y A VDD VDD pmos1v w=0.36u l=0.1u
.ends INVXL

* Spice subcircuit definition for MDFFHQX1




.subckt MDFFHQX1 Q / CK D0 D1 S0
mn10 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D0 VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 S0b D0b VSS nmos1v w=0.43u l=0.1u
mn13 n12 D1 VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 S0 D0b VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 D0b CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mp10 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D0 VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 S0 D0b VDD pmos1v w=0.65u l=0.1u
mp13 n13 D1 VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 S0b D0b VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 D0b CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
.ends MDFFHQX1

* Spice subcircuit definition for MDFFHQX2




.subckt MDFFHQX2 Q / CK D0 D1 S0
mn10 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D0 VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 S0b D0b VSS nmos1v w=0.43u l=0.1u
mn13 n12 D1 VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 S0 D0b VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 D0b CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mp10 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D0 VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 S0 D0b VDD pmos1v w=0.65u l=0.1u
mp13 n13 D1 VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 S0b D0b VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 D0b CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
.ends MDFFHQX2

* Spice subcircuit definition for MDFFHQX4




.subckt MDFFHQX4 Q / CK D0 D1 S0
mn10 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D0 VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 S0b D0b VSS nmos1v w=0.43u l=0.1u
mn13 n12 D1 VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 S0 D0b VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 D0b CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mp10 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D0 VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 S0 D0b VDD pmos1v w=0.65u l=0.1u
mp13 n13 D1 VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 S0b D0b VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 D0b CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
.ends MDFFHQX4

* Spice subcircuit definition for MDFFHQX8




.subckt MDFFHQX8 Q / CK D0 D1 S0
mn10 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D0 VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 S0b D0b VSS nmos1v w=0.43u l=0.1u
mn13 n12 D1 VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 S0 D0b VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 D0b CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=1.29u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=3.44u l=0.1u
mp10 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D0 VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 S0 D0b VDD pmos1v w=0.65u l=0.1u
mp13 n13 D1 VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 S0b D0b VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 D0b CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.95u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=5.2u l=0.1u
.ends MDFFHQX8

* Spice subcircuit definition for MX2X1




.subckt MX2X1 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends MX2X1

* Spice subcircuit definition for MX2X2




.subckt MX2X2 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends MX2X2

* Spice subcircuit definition for MX2X4




.subckt MX2X4 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.34u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.34u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.34u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.34u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.52u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.52u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.52u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.52u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends MX2X4

* Spice subcircuit definition for MX2X6




.subckt MX2X6 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.34u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.34u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.34u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.34u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=2.58u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.52u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.52u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.52u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.52u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=3.9u l=0.1u
.ends MX2X6

* Spice subcircuit definition for MX2X8




.subckt MX2X8 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.34u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.34u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.34u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.34u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=3.44u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.52u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.52u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.52u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.52u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=5.2u l=0.1u
.ends MX2X8

* Spice subcircuit definition for MX2XL




.subckt MX2XL Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
.ends MX2XL

* Spice subcircuit definition for MX3X1




.subckt MX3X1 Y / A B C S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n4 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n4 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 n0 S1b n1 VSS nmos1v w=0.24u l=0.1u
mn7 n6 C VSS VSS nmos1v w=0.24u l=0.1u
mn8 n6 S1 n1 VSS nmos1v w=0.24u l=0.1u
mn9 Y n1 VSS VSS nmos1v w=0.43u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n5 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n5 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 n0 S1 n1 VDD pmos1v w=0.36u l=0.1u
mp7 n7 C VDD VDD pmos1v w=0.36u l=0.1u
mp8 n7 S1b n1 VDD pmos1v w=0.36u l=0.1u
mp9 Y n1 VDD VDD pmos1v w=0.65u l=0.1u
.ends MX3X1

* Spice subcircuit definition for MX3X2




.subckt MX3X2 Y / A B C S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n4 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n4 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 n0 S1b n1 VSS nmos1v w=0.24u l=0.1u
mn7 n6 C VSS VSS nmos1v w=0.24u l=0.1u
mn8 n6 S1 n1 VSS nmos1v w=0.24u l=0.1u
mn9 Y n1 VSS VSS nmos1v w=0.86u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n5 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n5 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 n0 S1 n1 VDD pmos1v w=0.36u l=0.1u
mp7 n7 C VDD VDD pmos1v w=0.36u l=0.1u
mp8 n7 S1b n1 VDD pmos1v w=0.36u l=0.1u
mp9 Y n1 VDD VDD pmos1v w=1.3u l=0.1u
.ends MX3X2

* Spice subcircuit definition for MX3X4




.subckt MX3X4 Y / A B C S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n4 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n4 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 n0 S1b n1 VSS nmos1v w=0.43u l=0.1u
mn7 n6 C VSS VSS nmos1v w=0.43u l=0.1u
mn8 n6 S1 n1 VSS nmos1v w=0.43u l=0.1u
mn9 Y n1 VSS VSS nmos1v w=1.72u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n5 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n5 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 n0 S1 n1 VDD pmos1v w=0.65u l=0.1u
mp7 n7 C VDD VDD pmos1v w=0.65u l=0.1u
mp8 n7 S1b n1 VDD pmos1v w=0.65u l=0.1u
mp9 Y n1 VDD VDD pmos1v w=2.6u l=0.1u
.ends MX3X4

* Spice subcircuit definition for MX3XL




.subckt MX3XL Y / A B C S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n4 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n4 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 n0 S1b n1 VSS nmos1v w=0.24u l=0.1u
mn7 n6 C VSS VSS nmos1v w=0.24u l=0.1u
mn8 n6 S1 n1 VSS nmos1v w=0.24u l=0.1u
mn9 Y n1 VSS VSS nmos1v w=0.24u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n5 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n5 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 n0 S1 n1 VDD pmos1v w=0.36u l=0.1u
mp7 n7 C VDD VDD pmos1v w=0.36u l=0.1u
mp8 n7 S1b n1 VDD pmos1v w=0.36u l=0.1u
mp9 Y n1 VDD VDD pmos1v w=0.36u l=0.1u
.ends MX3XL

* Spice subcircuit definition for MX4X1




.subckt MX4X1 Y / A B C D S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n0 S1b n2 VSS nmos1v w=0.24u l=0.1u
mn11 n1 S1 n2 VSS nmos1v w=0.24u l=0.1u
mn12 Y n2 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 n7 C VSS VSS nmos1v w=0.24u l=0.1u
mn7 n7 S0b n1 VSS nmos1v w=0.24u l=0.1u
mn8 n9 D VSS VSS nmos1v w=0.24u l=0.1u
mn9 n9 S0 n1 VSS nmos1v w=0.24u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n0 S1 n2 VDD pmos1v w=0.36u l=0.1u
mp11 n1 S1b n2 VDD pmos1v w=0.36u l=0.1u
mp12 Y n2 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 n8 C VDD VDD pmos1v w=0.36u l=0.1u
mp7 n8 S0 n1 VDD pmos1v w=0.36u l=0.1u
mp8 n10 D VDD VDD pmos1v w=0.36u l=0.1u
mp9 n10 S0b n1 VDD pmos1v w=0.36u l=0.1u
.ends MX4X1

* Spice subcircuit definition for MX4X2




.subckt MX4X2 Y / A B C D S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n0 S1b n2 VSS nmos1v w=0.24u l=0.1u
mn11 n1 S1 n2 VSS nmos1v w=0.24u l=0.1u
mn12 Y n2 VSS VSS nmos1v w=0.86u l=0.1u
mn2 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 n7 C VSS VSS nmos1v w=0.24u l=0.1u
mn7 n7 S0b n1 VSS nmos1v w=0.24u l=0.1u
mn8 n9 D VSS VSS nmos1v w=0.24u l=0.1u
mn9 n9 S0 n1 VSS nmos1v w=0.24u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n0 S1 n2 VDD pmos1v w=0.36u l=0.1u
mp11 n1 S1b n2 VDD pmos1v w=0.36u l=0.1u
mp12 Y n2 VDD VDD pmos1v w=1.3u l=0.1u
mp2 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 n8 C VDD VDD pmos1v w=0.36u l=0.1u
mp7 n8 S0 n1 VDD pmos1v w=0.36u l=0.1u
mp8 n10 D VDD VDD pmos1v w=0.36u l=0.1u
mp9 n10 S0b n1 VDD pmos1v w=0.36u l=0.1u
.ends MX4X2

* Spice subcircuit definition for MX4X4




.subckt MX4X4 Y / A B C D S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n0 S1b n2 VSS nmos1v w=0.43u l=0.1u
mn11 n1 S1 n2 VSS nmos1v w=0.43u l=0.1u
mn12 Y n2 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 n7 C VSS VSS nmos1v w=0.24u l=0.1u
mn7 n7 S0b n1 VSS nmos1v w=0.24u l=0.1u
mn8 n9 D VSS VSS nmos1v w=0.24u l=0.1u
mn9 n9 S0 n1 VSS nmos1v w=0.24u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n0 S1 n2 VDD pmos1v w=0.65u l=0.1u
mp11 n1 S1b n2 VDD pmos1v w=0.65u l=0.1u
mp12 Y n2 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 n8 C VDD VDD pmos1v w=0.36u l=0.1u
mp7 n8 S0 n1 VDD pmos1v w=0.36u l=0.1u
mp8 n10 D VDD VDD pmos1v w=0.36u l=0.1u
mp9 n10 S0b n1 VDD pmos1v w=0.36u l=0.1u
.ends MX4X4

* Spice subcircuit definition for MX4XL




.subckt MX4XL Y / A B C D S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n0 S1b n2 VSS nmos1v w=0.24u l=0.1u
mn11 n1 S1 n2 VSS nmos1v w=0.24u l=0.1u
mn12 Y n2 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 n7 C VSS VSS nmos1v w=0.24u l=0.1u
mn7 n7 S0b n1 VSS nmos1v w=0.24u l=0.1u
mn8 n9 D VSS VSS nmos1v w=0.24u l=0.1u
mn9 n9 S0 n1 VSS nmos1v w=0.24u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n0 S1 n2 VDD pmos1v w=0.36u l=0.1u
mp11 n1 S1b n2 VDD pmos1v w=0.36u l=0.1u
mp12 Y n2 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 n8 C VDD VDD pmos1v w=0.36u l=0.1u
mp7 n8 S0 n1 VDD pmos1v w=0.36u l=0.1u
mp8 n10 D VDD VDD pmos1v w=0.36u l=0.1u
mp9 n10 S0b n1 VDD pmos1v w=0.36u l=0.1u
.ends MX4XL

* Spice subcircuit definition for MXI2X1




.subckt MXI2X1 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.43u l=0.1u
mn2 n3 S0b Y VSS nmos1v w=0.43u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.43u l=0.1u
mn4 n5 S0 Y VSS nmos1v w=0.43u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.65u l=0.1u
mp2 n4 S0 Y VDD pmos1v w=0.65u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.65u l=0.1u
mp4 n6 S0b Y VDD pmos1v w=0.65u l=0.1u
.ends MXI2X1

* Spice subcircuit definition for MXI2X2




.subckt MXI2X2 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn5 n1 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn6 Y n1 VSS VSS nmos1v w=0.86u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp5 n1 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp6 Y n1 VDD VDD pmos1v w=1.3u l=0.1u
.ends MXI2X2

* Spice subcircuit definition for MXI2X4




.subckt MXI2X4 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn5 n1 n0 VSS VSS nmos1v w=0.43u l=0.1u
mn6 Y n1 VSS VSS nmos1v w=1.72u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp5 n1 n0 VDD VDD pmos1v w=0.65u l=0.1u
mp6 Y n1 VDD VDD pmos1v w=2.6u l=0.1u
.ends MXI2X4

* Spice subcircuit definition for MXI2X6




.subckt MXI2X6 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn5 n1 n0 VSS VSS nmos1v w=0.86u l=0.1u
mn6 Y n1 VSS VSS nmos1v w=2.58u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp5 n1 n0 VDD VDD pmos1v w=1.3u l=0.1u
mp6 Y n1 VDD VDD pmos1v w=3.9u l=0.1u
.ends MXI2X6

* Spice subcircuit definition for MXI2X8




.subckt MXI2X8 Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn4 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn5 n1 n0 VSS VSS nmos1v w=0.86u l=0.1u
mn6 Y n1 VSS VSS nmos1v w=3.44u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp4 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp5 n1 n0 VDD VDD pmos1v w=1.3u l=0.1u
mp6 Y n1 VDD VDD pmos1v w=5.2u l=0.1u
.ends MXI2X8

* Spice subcircuit definition for MXI2XL




.subckt MXI2XL Y / A B S0
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 S0b Y VSS nmos1v w=0.24u l=0.1u
mn3 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn4 n5 S0 Y VSS nmos1v w=0.24u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 S0 Y VDD pmos1v w=0.36u l=0.1u
mp3 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp4 n6 S0b Y VDD pmos1v w=0.36u l=0.1u
.ends MXI2XL

* Spice subcircuit definition for MXI3X1




.subckt MXI3X1 Y / A B C S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n8 S1 n1 VSS nmos1v w=0.24u l=0.1u
mn11 Y n1 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n4 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n4 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 Cp C VSS VSS nmos1v w=0.24u l=0.1u
mn7 n6 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn8 n6 S1b n1 VSS nmos1v w=0.24u l=0.1u
mn9 n8 Cp VSS VSS nmos1v w=0.24u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n9 S1b n1 VDD pmos1v w=0.36u l=0.1u
mp11 Y n1 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n5 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n5 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 Cp C VDD VDD pmos1v w=0.36u l=0.1u
mp7 n7 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp8 n7 S1 n1 VDD pmos1v w=0.36u l=0.1u
mp9 n9 Cp VDD VDD pmos1v w=0.36u l=0.1u
.ends MXI3X1

* Spice subcircuit definition for MXI3X2




.subckt MXI3X2 Y / A B C S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n8 S1 n1 VSS nmos1v w=0.24u l=0.1u
mn11 Y n1 VSS VSS nmos1v w=0.86u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n4 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n4 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 Cp C VSS VSS nmos1v w=0.24u l=0.1u
mn7 n6 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn8 n6 S1b n1 VSS nmos1v w=0.24u l=0.1u
mn9 n8 Cp VSS VSS nmos1v w=0.24u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n9 S1b n1 VDD pmos1v w=0.36u l=0.1u
mp11 Y n1 VDD VDD pmos1v w=1.3u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n5 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n5 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 Cp C VDD VDD pmos1v w=0.36u l=0.1u
mp7 n7 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp8 n7 S1 n1 VDD pmos1v w=0.36u l=0.1u
mp9 n9 Cp VDD VDD pmos1v w=0.36u l=0.1u
.ends MXI3X2

* Spice subcircuit definition for MXI3X4




.subckt MXI3X4 Y / A B C S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n8 S1 n1 VSS nmos1v w=0.34u l=0.1u
mn11 Y n1 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n4 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n4 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 Cp C VSS VSS nmos1v w=0.24u l=0.1u
mn7 n6 n0 VSS VSS nmos1v w=0.34u l=0.1u
mn8 n6 S1b n1 VSS nmos1v w=0.34u l=0.1u
mn9 n8 Cp VSS VSS nmos1v w=0.34u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n9 S1b n1 VDD pmos1v w=0.52u l=0.1u
mp11 Y n1 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n5 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n5 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 Cp C VDD VDD pmos1v w=0.36u l=0.1u
mp7 n7 n0 VDD VDD pmos1v w=0.52u l=0.1u
mp8 n7 S1 n1 VDD pmos1v w=0.52u l=0.1u
mp9 n9 Cp VDD VDD pmos1v w=0.52u l=0.1u
.ends MXI3X4

* Spice subcircuit definition for MXI3XL




.subckt MXI3XL Y / A B C S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n8 S1 n1 VSS nmos1v w=0.24u l=0.1u
mn11 Y n1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n4 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n4 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 Cp C VSS VSS nmos1v w=0.24u l=0.1u
mn7 n6 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn8 n6 S1b n1 VSS nmos1v w=0.24u l=0.1u
mn9 n8 Cp VSS VSS nmos1v w=0.24u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n9 S1b n1 VDD pmos1v w=0.36u l=0.1u
mp11 Y n1 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n5 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n5 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 Cp C VDD VDD pmos1v w=0.36u l=0.1u
mp7 n7 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp8 n7 S1 n1 VDD pmos1v w=0.36u l=0.1u
mp9 n9 Cp VDD VDD pmos1v w=0.36u l=0.1u
.ends MXI3XL

* Spice subcircuit definition for MXI4X1




.subckt MXI4X1 Y / A B C D S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n11 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn11 n11 S1b n2 VSS nmos1v w=0.24u l=0.1u
mn12 n13 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn13 n13 S1 n2 VSS nmos1v w=0.24u l=0.1u
mn14 Y n2 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 n7 C VSS VSS nmos1v w=0.24u l=0.1u
mn7 n7 S0b n1 VSS nmos1v w=0.24u l=0.1u
mn8 n9 D VSS VSS nmos1v w=0.24u l=0.1u
mn9 n9 S0 n1 VSS nmos1v w=0.24u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n12 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp11 n12 S1 n2 VDD pmos1v w=0.36u l=0.1u
mp12 n14 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp13 n14 S1b n2 VDD pmos1v w=0.36u l=0.1u
mp14 Y n2 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 n8 C VDD VDD pmos1v w=0.36u l=0.1u
mp7 n8 S0 n1 VDD pmos1v w=0.36u l=0.1u
mp8 n10 D VDD VDD pmos1v w=0.36u l=0.1u
mp9 n10 S0b n1 VDD pmos1v w=0.36u l=0.1u
.ends MXI4X1

* Spice subcircuit definition for MXI4X2




.subckt MXI4X2 Y / A B C D S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n11 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn11 n11 S1b n2 VSS nmos1v w=0.24u l=0.1u
mn12 n13 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn13 n13 S1 n2 VSS nmos1v w=0.24u l=0.1u
mn14 Y n2 VSS VSS nmos1v w=0.86u l=0.1u
mn2 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 n7 C VSS VSS nmos1v w=0.24u l=0.1u
mn7 n7 S0b n1 VSS nmos1v w=0.24u l=0.1u
mn8 n9 D VSS VSS nmos1v w=0.24u l=0.1u
mn9 n9 S0 n1 VSS nmos1v w=0.24u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n12 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp11 n12 S1 n2 VDD pmos1v w=0.36u l=0.1u
mp12 n14 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp13 n14 S1b n2 VDD pmos1v w=0.36u l=0.1u
mp14 Y n2 VDD VDD pmos1v w=1.3u l=0.1u
mp2 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 n8 C VDD VDD pmos1v w=0.36u l=0.1u
mp7 n8 S0 n1 VDD pmos1v w=0.36u l=0.1u
mp8 n10 D VDD VDD pmos1v w=0.36u l=0.1u
mp9 n10 S0b n1 VDD pmos1v w=0.36u l=0.1u
.ends MXI4X2

* Spice subcircuit definition for MXI4X4




.subckt MXI4X4 Y / A B C D S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n11 n0 VSS VSS nmos1v w=0.34u l=0.1u
mn11 n11 S1b n2 VSS nmos1v w=0.34u l=0.1u
mn12 n13 n1 VSS VSS nmos1v w=0.34u l=0.1u
mn13 n13 S1 n2 VSS nmos1v w=0.34u l=0.1u
mn14 Y n2 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 n7 C VSS VSS nmos1v w=0.24u l=0.1u
mn7 n7 S0b n1 VSS nmos1v w=0.24u l=0.1u
mn8 n9 D VSS VSS nmos1v w=0.24u l=0.1u
mn9 n9 S0 n1 VSS nmos1v w=0.24u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n12 n0 VDD VDD pmos1v w=0.52u l=0.1u
mp11 n12 S1 n2 VDD pmos1v w=0.52u l=0.1u
mp12 n14 n1 VDD VDD pmos1v w=0.52u l=0.1u
mp13 n14 S1b n2 VDD pmos1v w=0.52u l=0.1u
mp14 Y n2 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 n8 C VDD VDD pmos1v w=0.36u l=0.1u
mp7 n8 S0 n1 VDD pmos1v w=0.36u l=0.1u
mp8 n10 D VDD VDD pmos1v w=0.36u l=0.1u
mp9 n10 S0b n1 VDD pmos1v w=0.36u l=0.1u
.ends MXI4X4

* Spice subcircuit definition for MXI4XL




.subckt MXI4XL Y / A B C D S0 S1
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 S1b S1 VSS VSS nmos1v w=0.24u l=0.1u
mn10 n11 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn11 n11 S1b n2 VSS nmos1v w=0.24u l=0.1u
mn12 n13 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn13 n13 S1 n2 VSS nmos1v w=0.24u l=0.1u
mn14 Y n2 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 A VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 S0b n0 VSS nmos1v w=0.24u l=0.1u
mn4 n5 B VSS VSS nmos1v w=0.24u l=0.1u
mn5 n5 S0 n0 VSS nmos1v w=0.24u l=0.1u
mn6 n7 C VSS VSS nmos1v w=0.24u l=0.1u
mn7 n7 S0b n1 VSS nmos1v w=0.24u l=0.1u
mn8 n9 D VSS VSS nmos1v w=0.24u l=0.1u
mn9 n9 S0 n1 VSS nmos1v w=0.24u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 S1b S1 VDD VDD pmos1v w=0.36u l=0.1u
mp10 n12 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp11 n12 S1 n2 VDD pmos1v w=0.36u l=0.1u
mp12 n14 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp13 n14 S1b n2 VDD pmos1v w=0.36u l=0.1u
mp14 Y n2 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 A VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 S0 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n6 B VDD VDD pmos1v w=0.36u l=0.1u
mp5 n6 S0b n0 VDD pmos1v w=0.36u l=0.1u
mp6 n8 C VDD VDD pmos1v w=0.36u l=0.1u
mp7 n8 S0 n1 VDD pmos1v w=0.36u l=0.1u
mp8 n10 D VDD VDD pmos1v w=0.36u l=0.1u
mp9 n10 S0b n1 VDD pmos1v w=0.36u l=0.1u
.ends MXI4XL

* Spice subcircuit definition for NAND2BX1




.subckt NAND2BX1 Y / AN B
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 n0 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n1 B Y VSS nmos1v w=0.43u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
mp2 Y B VDD VDD pmos1v w=0.65u l=0.1u
.ends NAND2BX1

* Spice subcircuit definition for NAND2BX2




.subckt NAND2BX2 Y / AN B
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 n0 VSS VSS nmos1v w=0.86u l=0.1u
mn2 n1 B Y VSS nmos1v w=0.86u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
mp2 Y B VDD VDD pmos1v w=1.3u l=0.1u
.ends NAND2BX2

* Spice subcircuit definition for NAND2BX4




.subckt NAND2BX4 Y / AN B
mn0 n0 AN VSS VSS nmos1v w=0.43u l=0.1u
mn1 n1 n0 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n1 B Y VSS nmos1v w=1.72u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.65u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
mp2 Y B VDD VDD pmos1v w=2.6u l=0.1u
.ends NAND2BX4

* Spice subcircuit definition for NAND2BXL




.subckt NAND2BXL Y / AN B
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n1 B Y VSS nmos1v w=0.24u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
mp2 Y B VDD VDD pmos1v w=0.36u l=0.1u
.ends NAND2BXL

* Spice subcircuit definition for NAND2X1




.subckt NAND2X1 Y / A B
mn0 n0 A VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 B Y VSS nmos1v w=0.43u l=0.1u
mp0 Y A VDD VDD pmos1v w=0.65u l=0.1u
mp1 Y B VDD VDD pmos1v w=0.65u l=0.1u
.ends NAND2X1

* Spice subcircuit definition for NAND2X2




.subckt NAND2X2 Y / A B
mn0 n0 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 B Y VSS nmos1v w=0.86u l=0.1u
mp0 Y A VDD VDD pmos1v w=1.3u l=0.1u
mp1 Y B VDD VDD pmos1v w=1.3u l=0.1u
.ends NAND2X2

* Spice subcircuit definition for NAND2X4




.subckt NAND2X4 Y / A B
mn0 n0 A VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 B Y VSS nmos1v w=1.72u l=0.1u
mp0 Y A VDD VDD pmos1v w=2.6u l=0.1u
mp1 Y B VDD VDD pmos1v w=2.6u l=0.1u
.ends NAND2X4

* Spice subcircuit definition for NAND2X6




.subckt NAND2X6 Y / A B
mn0 n0 A VSS VSS nmos1v w=2.58u l=0.1u
mn1 n0 B Y VSS nmos1v w=2.58u l=0.1u
mp0 Y A VDD VDD pmos1v w=3.9u l=0.1u
mp1 Y B VDD VDD pmos1v w=3.9u l=0.1u
.ends NAND2X6

* Spice subcircuit definition for NAND2X8




.subckt NAND2X8 Y / A B
mn0 n0 A VSS VSS nmos1v w=3.44u l=0.1u
mn1 n0 B Y VSS nmos1v w=3.44u l=0.1u
mp0 Y A VDD VDD pmos1v w=5.2u l=0.1u
mp1 Y B VDD VDD pmos1v w=5.2u l=0.1u
.ends NAND2X8

* Spice subcircuit definition for NAND2XL




.subckt NAND2XL Y / A B
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 B Y VSS nmos1v w=0.24u l=0.1u
mp0 Y A VDD VDD pmos1v w=0.36u l=0.1u
mp1 Y B VDD VDD pmos1v w=0.36u l=0.1u
.ends NAND2XL

* Spice subcircuit definition for NAND3BX1




.subckt NAND3BX1 Y / AN B C
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 n0 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n1 B n2 VSS nmos1v w=0.43u l=0.1u
mn3 n2 C Y VSS nmos1v w=0.43u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
mp2 Y B VDD VDD pmos1v w=0.65u l=0.1u
mp3 Y C VDD VDD pmos1v w=0.65u l=0.1u
.ends NAND3BX1

* Spice subcircuit definition for NAND3BX2




.subckt NAND3BX2 Y / AN B C
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 n0 VSS VSS nmos1v w=0.86u l=0.1u
mn2 n1 B n2 VSS nmos1v w=0.86u l=0.1u
mn3 n2 C Y VSS nmos1v w=0.86u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
mp2 Y B VDD VDD pmos1v w=1.3u l=0.1u
mp3 Y C VDD VDD pmos1v w=1.3u l=0.1u
.ends NAND3BX2

* Spice subcircuit definition for NAND3BX4




.subckt NAND3BX4 Y / AN B C
mn0 n0 AN VSS VSS nmos1v w=0.43u l=0.1u
mn1 n1 n0 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n1 B n2 VSS nmos1v w=1.72u l=0.1u
mn3 n2 C Y VSS nmos1v w=1.72u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.65u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
mp2 Y B VDD VDD pmos1v w=2.6u l=0.1u
mp3 Y C VDD VDD pmos1v w=2.6u l=0.1u
.ends NAND3BX4

* Spice subcircuit definition for NAND3BXL




.subckt NAND3BXL Y / AN B C
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n1 B n2 VSS nmos1v w=0.24u l=0.1u
mn3 n2 C Y VSS nmos1v w=0.24u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
mp2 Y B VDD VDD pmos1v w=0.36u l=0.1u
mp3 Y C VDD VDD pmos1v w=0.36u l=0.1u
.ends NAND3BXL

* Spice subcircuit definition for NAND3X1




.subckt NAND3X1 Y / A B C
mn0 n0 A VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 B n1 VSS nmos1v w=0.43u l=0.1u
mn2 n1 C Y VSS nmos1v w=0.43u l=0.1u
mp0 Y A VDD VDD pmos1v w=0.65u l=0.1u
mp1 Y B VDD VDD pmos1v w=0.65u l=0.1u
mp2 Y C VDD VDD pmos1v w=0.65u l=0.1u
.ends NAND3X1

* Spice subcircuit definition for NAND3X2




.subckt NAND3X2 Y / A B C
mn0 n0 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 B n1 VSS nmos1v w=0.86u l=0.1u
mn2 n1 C Y VSS nmos1v w=0.86u l=0.1u
mp0 Y A VDD VDD pmos1v w=1.3u l=0.1u
mp1 Y B VDD VDD pmos1v w=1.3u l=0.1u
mp2 Y C VDD VDD pmos1v w=1.3u l=0.1u
.ends NAND3X2

* Spice subcircuit definition for NAND3X4




.subckt NAND3X4 Y / A B C
mn0 n0 A VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 B n1 VSS nmos1v w=1.72u l=0.1u
mn2 n1 C Y VSS nmos1v w=1.72u l=0.1u
mp0 Y A VDD VDD pmos1v w=2.6u l=0.1u
mp1 Y B VDD VDD pmos1v w=2.6u l=0.1u
mp2 Y C VDD VDD pmos1v w=2.6u l=0.1u
.ends NAND3X4

* Spice subcircuit definition for NAND3X6




.subckt NAND3X6 Y / A B C
mn0 n0 A VSS VSS nmos1v w=2.58u l=0.1u
mn1 n0 B n1 VSS nmos1v w=2.58u l=0.1u
mn2 n1 C Y VSS nmos1v w=2.58u l=0.1u
mp0 Y A VDD VDD pmos1v w=3.9u l=0.1u
mp1 Y B VDD VDD pmos1v w=3.9u l=0.1u
mp2 Y C VDD VDD pmos1v w=3.9u l=0.1u
.ends NAND3X6

* Spice subcircuit definition for NAND3X8




.subckt NAND3X8 Y / A B C
mn0 n0 A VSS VSS nmos1v w=3.44u l=0.1u
mn1 n0 B n1 VSS nmos1v w=3.44u l=0.1u
mn2 n1 C Y VSS nmos1v w=3.44u l=0.1u
mp0 Y A VDD VDD pmos1v w=5.2u l=0.1u
mp1 Y B VDD VDD pmos1v w=5.2u l=0.1u
mp2 Y C VDD VDD pmos1v w=5.2u l=0.1u
.ends NAND3X8

* Spice subcircuit definition for NAND3XL




.subckt NAND3XL Y / A B C
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 B n1 VSS nmos1v w=0.24u l=0.1u
mn2 n1 C Y VSS nmos1v w=0.24u l=0.1u
mp0 Y A VDD VDD pmos1v w=0.36u l=0.1u
mp1 Y B VDD VDD pmos1v w=0.36u l=0.1u
mp2 Y C VDD VDD pmos1v w=0.36u l=0.1u
.ends NAND3XL

* Spice subcircuit definition for NAND4BBX1




.subckt NAND4BBX1 Y / AN BN C D
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 BN VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=0.43u l=0.1u
mn3 n2 n1 n3 VSS nmos1v w=0.43u l=0.1u
mn4 n3 C n4 VSS nmos1v w=0.43u l=0.1u
mn5 n4 D Y VSS nmos1v w=0.43u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 BN VDD VDD pmos1v w=0.36u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
mp3 Y n1 VDD VDD pmos1v w=0.65u l=0.1u
mp4 Y C VDD VDD pmos1v w=0.65u l=0.1u
mp5 Y D VDD VDD pmos1v w=0.65u l=0.1u
.ends NAND4BBX1

* Spice subcircuit definition for NAND4BBX2




.subckt NAND4BBX2 Y / AN BN C D
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 BN VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=0.86u l=0.1u
mn3 n2 n1 n3 VSS nmos1v w=0.86u l=0.1u
mn4 n3 C n4 VSS nmos1v w=0.86u l=0.1u
mn5 n4 D Y VSS nmos1v w=0.86u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 BN VDD VDD pmos1v w=0.36u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
mp3 Y n1 VDD VDD pmos1v w=1.3u l=0.1u
mp4 Y C VDD VDD pmos1v w=1.3u l=0.1u
mp5 Y D VDD VDD pmos1v w=1.3u l=0.1u
.ends NAND4BBX2

* Spice subcircuit definition for NAND4BBX4




.subckt NAND4BBX4 Y / AN BN C D
mn0 n0 AN VSS VSS nmos1v w=0.43u l=0.1u
mn1 n1 BN VSS VSS nmos1v w=0.43u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=1.72u l=0.1u
mn3 n2 n1 n3 VSS nmos1v w=1.72u l=0.1u
mn4 n3 C n4 VSS nmos1v w=1.72u l=0.1u
mn5 n4 D Y VSS nmos1v w=1.72u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 BN VDD VDD pmos1v w=0.65u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
mp3 Y n1 VDD VDD pmos1v w=2.6u l=0.1u
mp4 Y C VDD VDD pmos1v w=2.6u l=0.1u
mp5 Y D VDD VDD pmos1v w=2.6u l=0.1u
.ends NAND4BBX4

* Spice subcircuit definition for NAND4BBXL




.subckt NAND4BBXL Y / AN BN C D
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 BN VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 n1 n3 VSS nmos1v w=0.24u l=0.1u
mn4 n3 C n4 VSS nmos1v w=0.24u l=0.1u
mn5 n4 D Y VSS nmos1v w=0.24u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 BN VDD VDD pmos1v w=0.36u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 Y n1 VDD VDD pmos1v w=0.36u l=0.1u
mp4 Y C VDD VDD pmos1v w=0.36u l=0.1u
mp5 Y D VDD VDD pmos1v w=0.36u l=0.1u
.ends NAND4BBXL

* Spice subcircuit definition for NAND4BX1




.subckt NAND4BX1 Y / AN B C D
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 n0 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n1 B n2 VSS nmos1v w=0.43u l=0.1u
mn3 n2 C n3 VSS nmos1v w=0.43u l=0.1u
mn4 n3 D Y VSS nmos1v w=0.43u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
mp2 Y B VDD VDD pmos1v w=0.65u l=0.1u
mp3 Y C VDD VDD pmos1v w=0.65u l=0.1u
mp4 Y D VDD VDD pmos1v w=0.65u l=0.1u
.ends NAND4BX1

* Spice subcircuit definition for NAND4BX2




.subckt NAND4BX2 Y / AN B C D
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 n0 VSS VSS nmos1v w=0.86u l=0.1u
mn2 n1 B n2 VSS nmos1v w=0.86u l=0.1u
mn3 n2 C n3 VSS nmos1v w=0.86u l=0.1u
mn4 n3 D Y VSS nmos1v w=0.86u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
mp2 Y B VDD VDD pmos1v w=1.3u l=0.1u
mp3 Y C VDD VDD pmos1v w=1.3u l=0.1u
mp4 Y D VDD VDD pmos1v w=1.3u l=0.1u
.ends NAND4BX2

* Spice subcircuit definition for NAND4BX4




.subckt NAND4BX4 Y / AN B C D
mn0 n0 AN VSS VSS nmos1v w=0.43u l=0.1u
mn1 n1 n0 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n1 B n2 VSS nmos1v w=1.72u l=0.1u
mn3 n2 C n3 VSS nmos1v w=1.72u l=0.1u
mn4 n3 D Y VSS nmos1v w=1.72u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.65u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
mp2 Y B VDD VDD pmos1v w=2.6u l=0.1u
mp3 Y C VDD VDD pmos1v w=2.6u l=0.1u
mp4 Y D VDD VDD pmos1v w=2.6u l=0.1u
.ends NAND4BX4

* Spice subcircuit definition for NAND4BXL




.subckt NAND4BXL Y / AN B C D
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n1 B n2 VSS nmos1v w=0.24u l=0.1u
mn3 n2 C n3 VSS nmos1v w=0.24u l=0.1u
mn4 n3 D Y VSS nmos1v w=0.24u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
mp2 Y B VDD VDD pmos1v w=0.36u l=0.1u
mp3 Y C VDD VDD pmos1v w=0.36u l=0.1u
mp4 Y D VDD VDD pmos1v w=0.36u l=0.1u
.ends NAND4BXL

* Spice subcircuit definition for NAND4X1




.subckt NAND4X1 Y / A B C D
mn0 n0 A VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 B n1 VSS nmos1v w=0.43u l=0.1u
mn2 n1 C n2 VSS nmos1v w=0.43u l=0.1u
mn3 n2 D Y VSS nmos1v w=0.43u l=0.1u
mp0 Y A VDD VDD pmos1v w=0.65u l=0.1u
mp1 Y B VDD VDD pmos1v w=0.65u l=0.1u
mp2 Y C VDD VDD pmos1v w=0.65u l=0.1u
mp3 Y D VDD VDD pmos1v w=0.65u l=0.1u
.ends NAND4X1

* Spice subcircuit definition for NAND4X2




.subckt NAND4X2 Y / A B C D
mn0 n0 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 B n1 VSS nmos1v w=0.86u l=0.1u
mn2 n1 C n2 VSS nmos1v w=0.86u l=0.1u
mn3 n2 D Y VSS nmos1v w=0.86u l=0.1u
mp0 Y A VDD VDD pmos1v w=1.3u l=0.1u
mp1 Y B VDD VDD pmos1v w=1.3u l=0.1u
mp2 Y C VDD VDD pmos1v w=1.3u l=0.1u
mp3 Y D VDD VDD pmos1v w=1.3u l=0.1u
.ends NAND4X2

* Spice subcircuit definition for NAND4X4




.subckt NAND4X4 Y / A B C D
mn0 n0 A VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 B n1 VSS nmos1v w=1.72u l=0.1u
mn2 n1 C n2 VSS nmos1v w=1.72u l=0.1u
mn3 n2 D Y VSS nmos1v w=1.72u l=0.1u
mp0 Y A VDD VDD pmos1v w=2.6u l=0.1u
mp1 Y B VDD VDD pmos1v w=2.6u l=0.1u
mp2 Y C VDD VDD pmos1v w=2.6u l=0.1u
mp3 Y D VDD VDD pmos1v w=2.6u l=0.1u
.ends NAND4X4

* Spice subcircuit definition for NAND4X6




.subckt NAND4X6 Y / A B C D
mn0 n0 A VSS VSS nmos1v w=2.58u l=0.1u
mn1 n0 B n1 VSS nmos1v w=2.58u l=0.1u
mn2 n1 C n2 VSS nmos1v w=2.58u l=0.1u
mn3 n2 D Y VSS nmos1v w=2.58u l=0.1u
mp0 Y A VDD VDD pmos1v w=3.9u l=0.1u
mp1 Y B VDD VDD pmos1v w=3.9u l=0.1u
mp2 Y C VDD VDD pmos1v w=3.9u l=0.1u
mp3 Y D VDD VDD pmos1v w=3.9u l=0.1u
.ends NAND4X6

* Spice subcircuit definition for NAND4X8




.subckt NAND4X8 Y / A B C D
mn0 n0 A VSS VSS nmos1v w=3.44u l=0.1u
mn1 n0 B n1 VSS nmos1v w=3.44u l=0.1u
mn2 n1 C n2 VSS nmos1v w=3.44u l=0.1u
mn3 n2 D Y VSS nmos1v w=3.44u l=0.1u
mp0 Y A VDD VDD pmos1v w=5.2u l=0.1u
mp1 Y B VDD VDD pmos1v w=5.2u l=0.1u
mp2 Y C VDD VDD pmos1v w=5.2u l=0.1u
mp3 Y D VDD VDD pmos1v w=5.2u l=0.1u
.ends NAND4X8

* Spice subcircuit definition for NAND4XL




.subckt NAND4XL Y / A B C D
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 B n1 VSS nmos1v w=0.24u l=0.1u
mn2 n1 C n2 VSS nmos1v w=0.24u l=0.1u
mn3 n2 D Y VSS nmos1v w=0.24u l=0.1u
mp0 Y A VDD VDD pmos1v w=0.36u l=0.1u
mp1 Y B VDD VDD pmos1v w=0.36u l=0.1u
mp2 Y C VDD VDD pmos1v w=0.36u l=0.1u
mp3 Y D VDD VDD pmos1v w=0.36u l=0.1u
.ends NAND4XL

* Spice subcircuit definition for NOR2BX1




.subckt NOR2BX1 Y / AN B
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mn2 Y B VSS VSS nmos1v w=0.43u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 n0 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n1 B Y VDD pmos1v w=0.65u l=0.1u
.ends NOR2BX1

* Spice subcircuit definition for NOR2BX2




.subckt NOR2BX2 Y / AN B
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mn2 Y B VSS VSS nmos1v w=0.86u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 n0 VDD VDD pmos1v w=1.3u l=0.1u
mp2 n1 B Y VDD pmos1v w=1.3u l=0.1u
.ends NOR2BX2

* Spice subcircuit definition for NOR2BX4




.subckt NOR2BX4 Y / AN B
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mn2 Y B VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 n0 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n1 B Y VDD pmos1v w=2.6u l=0.1u
.ends NOR2BX4

* Spice subcircuit definition for NOR2BXL




.subckt NOR2BXL Y / AN B
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mn2 Y B VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n1 B Y VDD pmos1v w=0.36u l=0.1u
.ends NOR2BXL

* Spice subcircuit definition for NOR2X1




.subckt NOR2X1 Y / A B
mn0 Y A VSS VSS nmos1v w=0.43u l=0.1u
mn1 Y B VSS VSS nmos1v w=0.43u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 n0 B Y VDD pmos1v w=0.65u l=0.1u
.ends NOR2X1

* Spice subcircuit definition for NOR2X2




.subckt NOR2X2 Y / A B
mn0 Y A VSS VSS nmos1v w=0.86u l=0.1u
mn1 Y B VSS VSS nmos1v w=0.86u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n0 B Y VDD pmos1v w=1.3u l=0.1u
.ends NOR2X2

* Spice subcircuit definition for NOR2X4




.subckt NOR2X4 Y / A B
mn0 Y A VSS VSS nmos1v w=1.72u l=0.1u
mn1 Y B VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 A VDD VDD pmos1v w=2.6u l=0.1u
mp1 n0 B Y VDD pmos1v w=2.6u l=0.1u
.ends NOR2X4

* Spice subcircuit definition for NOR2X6




.subckt NOR2X6 Y / A B
mn0 Y A VSS VSS nmos1v w=2.58u l=0.1u
mn1 Y B VSS VSS nmos1v w=2.58u l=0.1u
mp0 n0 A VDD VDD pmos1v w=3.9u l=0.1u
mp1 n0 B Y VDD pmos1v w=3.9u l=0.1u
.ends NOR2X6

* Spice subcircuit definition for NOR2X8




.subckt NOR2X8 Y / A B
mn0 Y A VSS VSS nmos1v w=3.44u l=0.1u
mn1 Y B VSS VSS nmos1v w=3.44u l=0.1u
mp0 n0 A VDD VDD pmos1v w=5.2u l=0.1u
mp1 n0 B Y VDD pmos1v w=5.2u l=0.1u
.ends NOR2X8

* Spice subcircuit definition for NOR2XL




.subckt NOR2XL Y / A B
mn0 Y A VSS VSS nmos1v w=0.24u l=0.1u
mn1 Y B VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 B Y VDD pmos1v w=0.36u l=0.1u
.ends NOR2XL

* Spice subcircuit definition for NOR3BX1




.subckt NOR3BX1 Y / AN B C
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mn2 Y B VSS VSS nmos1v w=0.43u l=0.1u
mn3 Y C VSS VSS nmos1v w=0.43u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 n0 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n1 B n2 VDD pmos1v w=0.65u l=0.1u
mp3 n2 C Y VDD pmos1v w=0.65u l=0.1u
.ends NOR3BX1

* Spice subcircuit definition for NOR3BX2




.subckt NOR3BX2 Y / AN B C
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mn2 Y B VSS VSS nmos1v w=0.86u l=0.1u
mn3 Y C VSS VSS nmos1v w=0.86u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 n0 VDD VDD pmos1v w=1.3u l=0.1u
mp2 n1 B n2 VDD pmos1v w=1.3u l=0.1u
mp3 n2 C Y VDD pmos1v w=1.3u l=0.1u
.ends NOR3BX2

* Spice subcircuit definition for NOR3BX4




.subckt NOR3BX4 Y / AN B C
mn0 n0 AN VSS VSS nmos1v w=0.43u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mn2 Y B VSS VSS nmos1v w=1.72u l=0.1u
mn3 Y C VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 n0 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n1 B n2 VDD pmos1v w=2.6u l=0.1u
mp3 n2 C Y VDD pmos1v w=2.6u l=0.1u
.ends NOR3BX4

* Spice subcircuit definition for NOR3BXL




.subckt NOR3BXL Y / AN B C
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mn2 Y B VSS VSS nmos1v w=0.24u l=0.1u
mn3 Y C VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n1 B n2 VDD pmos1v w=0.36u l=0.1u
mp3 n2 C Y VDD pmos1v w=0.36u l=0.1u
.ends NOR3BXL

* Spice subcircuit definition for NOR3X1




.subckt NOR3X1 Y / A B C
mn0 Y A VSS VSS nmos1v w=0.43u l=0.1u
mn1 Y B VSS VSS nmos1v w=0.43u l=0.1u
mn2 Y C VSS VSS nmos1v w=0.43u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 n0 B n1 VDD pmos1v w=0.65u l=0.1u
mp2 n1 C Y VDD pmos1v w=0.65u l=0.1u
.ends NOR3X1

* Spice subcircuit definition for NOR3X2




.subckt NOR3X2 Y / A B C
mn0 Y A VSS VSS nmos1v w=0.86u l=0.1u
mn1 Y B VSS VSS nmos1v w=0.86u l=0.1u
mn2 Y C VSS VSS nmos1v w=0.86u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n0 B n1 VDD pmos1v w=1.3u l=0.1u
mp2 n1 C Y VDD pmos1v w=1.3u l=0.1u
.ends NOR3X2

* Spice subcircuit definition for NOR3X4




.subckt NOR3X4 Y / A B C
mn0 Y A VSS VSS nmos1v w=1.72u l=0.1u
mn1 Y B VSS VSS nmos1v w=1.72u l=0.1u
mn2 Y C VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 A VDD VDD pmos1v w=2.6u l=0.1u
mp1 n0 B n1 VDD pmos1v w=2.6u l=0.1u
mp2 n1 C Y VDD pmos1v w=2.6u l=0.1u
.ends NOR3X4

* Spice subcircuit definition for NOR3X6




.subckt NOR3X6 Y / A B C
mn0 Y A VSS VSS nmos1v w=2.58u l=0.1u
mn1 Y B VSS VSS nmos1v w=2.58u l=0.1u
mn2 Y C VSS VSS nmos1v w=2.58u l=0.1u
mp0 n0 A VDD VDD pmos1v w=3.9u l=0.1u
mp1 n0 B n1 VDD pmos1v w=3.9u l=0.1u
mp2 n1 C Y VDD pmos1v w=3.9u l=0.1u
.ends NOR3X6

* Spice subcircuit definition for NOR3X8




.subckt NOR3X8 Y / A B C
mn0 Y A VSS VSS nmos1v w=3.44u l=0.1u
mn1 Y B VSS VSS nmos1v w=3.44u l=0.1u
mn2 Y C VSS VSS nmos1v w=3.44u l=0.1u
mp0 n0 A VDD VDD pmos1v w=5.2u l=0.1u
mp1 n0 B n1 VDD pmos1v w=5.2u l=0.1u
mp2 n1 C Y VDD pmos1v w=5.2u l=0.1u
.ends NOR3X8

* Spice subcircuit definition for NOR3XL




.subckt NOR3XL Y / A B C
mn0 Y A VSS VSS nmos1v w=0.24u l=0.1u
mn1 Y B VSS VSS nmos1v w=0.24u l=0.1u
mn2 Y C VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 B n1 VDD pmos1v w=0.36u l=0.1u
mp2 n1 C Y VDD pmos1v w=0.36u l=0.1u
.ends NOR3XL

* Spice subcircuit definition for NOR4BBX1




.subckt NOR4BBX1 Y / AN BN C D
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 BN VSS VSS nmos1v w=0.24u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mn3 Y n1 VSS VSS nmos1v w=0.43u l=0.1u
mn4 Y C VSS VSS nmos1v w=0.43u l=0.1u
mn5 Y D VSS VSS nmos1v w=0.43u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 BN VDD VDD pmos1v w=0.36u l=0.1u
mp2 n2 n0 VDD VDD pmos1v w=0.65u l=0.1u
mp3 n2 n1 n3 VDD pmos1v w=0.65u l=0.1u
mp4 n3 C n4 VDD pmos1v w=0.65u l=0.1u
mp5 n4 D Y VDD pmos1v w=0.65u l=0.1u
.ends NOR4BBX1

* Spice subcircuit definition for NOR4BBX2




.subckt NOR4BBX2 Y / AN BN C D
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 BN VSS VSS nmos1v w=0.24u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mn3 Y n1 VSS VSS nmos1v w=0.86u l=0.1u
mn4 Y C VSS VSS nmos1v w=0.86u l=0.1u
mn5 Y D VSS VSS nmos1v w=0.86u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 BN VDD VDD pmos1v w=0.36u l=0.1u
mp2 n2 n0 VDD VDD pmos1v w=1.3u l=0.1u
mp3 n2 n1 n3 VDD pmos1v w=1.3u l=0.1u
mp4 n3 C n4 VDD pmos1v w=1.3u l=0.1u
mp5 n4 D Y VDD pmos1v w=1.3u l=0.1u
.ends NOR4BBX2

* Spice subcircuit definition for NOR4BBX4




.subckt NOR4BBX4 Y / AN BN C D
mn0 n0 AN VSS VSS nmos1v w=0.43u l=0.1u
mn1 n1 BN VSS VSS nmos1v w=0.43u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mn3 Y n1 VSS VSS nmos1v w=1.72u l=0.1u
mn4 Y C VSS VSS nmos1v w=1.72u l=0.1u
mn5 Y D VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 BN VDD VDD pmos1v w=0.65u l=0.1u
mp2 n2 n0 VDD VDD pmos1v w=2.6u l=0.1u
mp3 n2 n1 n3 VDD pmos1v w=2.6u l=0.1u
mp4 n3 C n4 VDD pmos1v w=2.6u l=0.1u
mp5 n4 D Y VDD pmos1v w=2.6u l=0.1u
.ends NOR4BBX4

* Spice subcircuit definition for NOR4BBXL




.subckt NOR4BBXL Y / AN BN C D
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 BN VSS VSS nmos1v w=0.24u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 Y n1 VSS VSS nmos1v w=0.24u l=0.1u
mn4 Y C VSS VSS nmos1v w=0.24u l=0.1u
mn5 Y D VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 BN VDD VDD pmos1v w=0.36u l=0.1u
mp2 n2 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n2 n1 n3 VDD pmos1v w=0.36u l=0.1u
mp4 n3 C n4 VDD pmos1v w=0.36u l=0.1u
mp5 n4 D Y VDD pmos1v w=0.36u l=0.1u
.ends NOR4BBXL

* Spice subcircuit definition for NOR4BX1




.subckt NOR4BX1 Y / AN B C D
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mn2 Y B VSS VSS nmos1v w=0.43u l=0.1u
mn3 Y C VSS VSS nmos1v w=0.43u l=0.1u
mn4 Y D VSS VSS nmos1v w=0.43u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 n0 VDD VDD pmos1v w=0.65u l=0.1u
mp2 n1 B n2 VDD pmos1v w=0.65u l=0.1u
mp3 n2 C n3 VDD pmos1v w=0.65u l=0.1u
mp4 n3 D Y VDD pmos1v w=0.65u l=0.1u
.ends NOR4BX1

* Spice subcircuit definition for NOR4BX2




.subckt NOR4BX2 Y / AN B C D
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mn2 Y B VSS VSS nmos1v w=0.86u l=0.1u
mn3 Y C VSS VSS nmos1v w=0.86u l=0.1u
mn4 Y D VSS VSS nmos1v w=0.86u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 n0 VDD VDD pmos1v w=1.3u l=0.1u
mp2 n1 B n2 VDD pmos1v w=1.3u l=0.1u
mp3 n2 C n3 VDD pmos1v w=1.3u l=0.1u
mp4 n3 D Y VDD pmos1v w=1.3u l=0.1u
.ends NOR4BX2

* Spice subcircuit definition for NOR4BX4




.subckt NOR4BX4 Y / AN B C D
mn0 n0 AN VSS VSS nmos1v w=0.43u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mn2 Y B VSS VSS nmos1v w=1.72u l=0.1u
mn3 Y C VSS VSS nmos1v w=1.72u l=0.1u
mn4 Y D VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 n0 VDD VDD pmos1v w=2.6u l=0.1u
mp2 n1 B n2 VDD pmos1v w=2.6u l=0.1u
mp3 n2 C n3 VDD pmos1v w=2.6u l=0.1u
mp4 n3 D Y VDD pmos1v w=2.6u l=0.1u
.ends NOR4BX4

* Spice subcircuit definition for NOR4BXL




.subckt NOR4BXL Y / AN B C D
mn0 n0 AN VSS VSS nmos1v w=0.24u l=0.1u
mn1 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mn2 Y B VSS VSS nmos1v w=0.24u l=0.1u
mn3 Y C VSS VSS nmos1v w=0.24u l=0.1u
mn4 Y D VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 AN VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp2 n1 B n2 VDD pmos1v w=0.36u l=0.1u
mp3 n2 C n3 VDD pmos1v w=0.36u l=0.1u
mp4 n3 D Y VDD pmos1v w=0.36u l=0.1u
.ends NOR4BXL

* Spice subcircuit definition for NOR4X1




.subckt NOR4X1 Y / A B C D
mn0 Y A VSS VSS nmos1v w=0.43u l=0.1u
mn1 Y B VSS VSS nmos1v w=0.43u l=0.1u
mn2 Y C VSS VSS nmos1v w=0.43u l=0.1u
mn3 Y D VSS VSS nmos1v w=0.43u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 n0 B n1 VDD pmos1v w=0.65u l=0.1u
mp2 n1 C n2 VDD pmos1v w=0.65u l=0.1u
mp3 n2 D Y VDD pmos1v w=0.65u l=0.1u
.ends NOR4X1

* Spice subcircuit definition for NOR4X2




.subckt NOR4X2 Y / A B C D
mn0 Y A VSS VSS nmos1v w=0.86u l=0.1u
mn1 Y B VSS VSS nmos1v w=0.86u l=0.1u
mn2 Y C VSS VSS nmos1v w=0.86u l=0.1u
mn3 Y D VSS VSS nmos1v w=0.86u l=0.1u
mp0 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n0 B n1 VDD pmos1v w=1.3u l=0.1u
mp2 n1 C n2 VDD pmos1v w=1.3u l=0.1u
mp3 n2 D Y VDD pmos1v w=1.3u l=0.1u
.ends NOR4X2

* Spice subcircuit definition for NOR4X4




.subckt NOR4X4 Y / A B C D
mn0 Y A VSS VSS nmos1v w=1.72u l=0.1u
mn1 Y B VSS VSS nmos1v w=1.72u l=0.1u
mn2 Y C VSS VSS nmos1v w=1.72u l=0.1u
mn3 Y D VSS VSS nmos1v w=1.72u l=0.1u
mp0 n0 A VDD VDD pmos1v w=2.6u l=0.1u
mp1 n0 B n1 VDD pmos1v w=2.6u l=0.1u
mp2 n1 C n2 VDD pmos1v w=2.6u l=0.1u
mp3 n2 D Y VDD pmos1v w=2.6u l=0.1u
.ends NOR4X4

* Spice subcircuit definition for NOR4X6




.subckt NOR4X6 Y / A B C D
mn0 Y A VSS VSS nmos1v w=2.58u l=0.1u
mn1 Y B VSS VSS nmos1v w=2.58u l=0.1u
mn2 Y C VSS VSS nmos1v w=2.58u l=0.1u
mn3 Y D VSS VSS nmos1v w=2.58u l=0.1u
mp0 n0 A VDD VDD pmos1v w=3.9u l=0.1u
mp1 n0 B n1 VDD pmos1v w=3.9u l=0.1u
mp2 n1 C n2 VDD pmos1v w=3.9u l=0.1u
mp3 n2 D Y VDD pmos1v w=3.9u l=0.1u
.ends NOR4X6

* Spice subcircuit definition for NOR4X8




.subckt NOR4X8 Y / A B C D
mn0 Y A VSS VSS nmos1v w=3.44u l=0.1u
mn1 Y B VSS VSS nmos1v w=3.44u l=0.1u
mn2 Y C VSS VSS nmos1v w=3.44u l=0.1u
mn3 Y D VSS VSS nmos1v w=3.44u l=0.1u
mp0 n0 A VDD VDD pmos1v w=5.2u l=0.1u
mp1 n0 B n1 VDD pmos1v w=5.2u l=0.1u
mp2 n1 C n2 VDD pmos1v w=5.2u l=0.1u
mp3 n2 D Y VDD pmos1v w=5.2u l=0.1u
.ends NOR4X8

* Spice subcircuit definition for NOR4XL




.subckt NOR4XL Y / A B C D
mn0 Y A VSS VSS nmos1v w=0.24u l=0.1u
mn1 Y B VSS VSS nmos1v w=0.24u l=0.1u
mn2 Y C VSS VSS nmos1v w=0.24u l=0.1u
mn3 Y D VSS VSS nmos1v w=0.24u l=0.1u
mp0 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 B n1 VDD pmos1v w=0.36u l=0.1u
mp2 n1 C n2 VDD pmos1v w=0.36u l=0.1u
mp3 n2 D Y VDD pmos1v w=0.36u l=0.1u
.ends NOR4XL

* Spice subcircuit definition for OA21X1




.subckt OA21X1 Y / A0 A1 B0
mn0 n1 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n1 B0 n0 VSS nmos1v w=0.24u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 A1 n0 VDD pmos1v w=0.36u l=0.1u
mp2 n0 B0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends OA21X1

* Spice subcircuit definition for OA21X2




.subckt OA21X2 Y / A0 A1 B0
mn0 n1 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n1 B0 n0 VSS nmos1v w=0.24u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 A1 n0 VDD pmos1v w=0.36u l=0.1u
mp2 n0 B0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends OA21X2

* Spice subcircuit definition for OA21X4




.subckt OA21X4 Y / A0 A1 B0
mn0 n1 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n1 A1 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n1 B0 n0 VSS nmos1v w=0.43u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n2 A1 n0 VDD pmos1v w=0.65u l=0.1u
mp2 n0 B0 VDD VDD pmos1v w=0.65u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends OA21X4

* Spice subcircuit definition for OA21XL




.subckt OA21XL Y / A0 A1 B0
mn0 n1 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n1 B0 n0 VSS nmos1v w=0.24u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 A1 n0 VDD pmos1v w=0.36u l=0.1u
mp2 n0 B0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
.ends OA21XL

* Spice subcircuit definition for OA22X1




.subckt OA22X1 Y / A0 A1 B0 B1
mn0 n1 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n1 B0 n0 VSS nmos1v w=0.24u l=0.1u
mn3 n1 B1 n0 VSS nmos1v w=0.24u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 A1 n0 VDD pmos1v w=0.36u l=0.1u
mp2 n3 B0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 B1 n0 VDD pmos1v w=0.36u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends OA22X1

* Spice subcircuit definition for OA22X2




.subckt OA22X2 Y / A0 A1 B0 B1
mn0 n1 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n1 B0 n0 VSS nmos1v w=0.24u l=0.1u
mn3 n1 B1 n0 VSS nmos1v w=0.24u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 A1 n0 VDD pmos1v w=0.36u l=0.1u
mp2 n3 B0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 B1 n0 VDD pmos1v w=0.36u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends OA22X2

* Spice subcircuit definition for OA22X4




.subckt OA22X4 Y / A0 A1 B0 B1
mn0 n1 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n1 A1 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n1 B0 n0 VSS nmos1v w=0.43u l=0.1u
mn3 n1 B1 n0 VSS nmos1v w=0.43u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n2 A1 n0 VDD pmos1v w=0.65u l=0.1u
mp2 n3 B0 VDD VDD pmos1v w=0.65u l=0.1u
mp3 n3 B1 n0 VDD pmos1v w=0.65u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends OA22X4

* Spice subcircuit definition for OA22XL




.subckt OA22XL Y / A0 A1 B0 B1
mn0 n1 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n1 B0 n0 VSS nmos1v w=0.24u l=0.1u
mn3 n1 B1 n0 VSS nmos1v w=0.24u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 A1 n0 VDD pmos1v w=0.36u l=0.1u
mp2 n3 B0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 B1 n0 VDD pmos1v w=0.36u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
.ends OA22XL

* Spice subcircuit definition for OAI211X1




.subckt OAI211X1 Y / A0 A1 B0 C0
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n0 B0 n1 VSS nmos1v w=0.43u l=0.1u
mn3 n1 C0 Y VSS nmos1v w=0.43u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n2 A1 Y VDD pmos1v w=0.65u l=0.1u
mp2 Y B0 VDD VDD pmos1v w=0.65u l=0.1u
mp3 Y C0 VDD VDD pmos1v w=0.65u l=0.1u
.ends OAI211X1

* Spice subcircuit definition for OAI211X2




.subckt OAI211X2 Y / A0 A1 B0 C0
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.86u l=0.1u
mn2 n0 B0 n1 VSS nmos1v w=0.86u l=0.1u
mn3 n1 C0 Y VSS nmos1v w=0.86u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n2 A1 Y VDD pmos1v w=1.3u l=0.1u
mp2 Y B0 VDD VDD pmos1v w=1.3u l=0.1u
mp3 Y C0 VDD VDD pmos1v w=1.3u l=0.1u
.ends OAI211X2

* Spice subcircuit definition for OAI211X4




.subckt OAI211X4 Y / A0 A1 B0 C0
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n0 B0 n1 VSS nmos1v w=1.72u l=0.1u
mn3 n1 C0 Y VSS nmos1v w=1.72u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n2 A1 Y VDD pmos1v w=2.6u l=0.1u
mp2 Y B0 VDD VDD pmos1v w=2.6u l=0.1u
mp3 Y C0 VDD VDD pmos1v w=2.6u l=0.1u
.ends OAI211X4

* Spice subcircuit definition for OAI211XL




.subckt OAI211XL Y / A0 A1 B0 C0
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n0 B0 n1 VSS nmos1v w=0.24u l=0.1u
mn3 n1 C0 Y VSS nmos1v w=0.24u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 A1 Y VDD pmos1v w=0.36u l=0.1u
mp2 Y B0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 Y C0 VDD VDD pmos1v w=0.36u l=0.1u
.ends OAI211XL

* Spice subcircuit definition for OAI21X1




.subckt OAI21X1 Y / A0 A1 B0
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n0 B0 Y VSS nmos1v w=0.43u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 A1 Y VDD pmos1v w=0.65u l=0.1u
mp2 Y B0 VDD VDD pmos1v w=0.65u l=0.1u
.ends OAI21X1

* Spice subcircuit definition for OAI21X2




.subckt OAI21X2 Y / A0 A1 B0
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.86u l=0.1u
mn2 n0 B0 Y VSS nmos1v w=0.86u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n1 A1 Y VDD pmos1v w=1.3u l=0.1u
mp2 Y B0 VDD VDD pmos1v w=1.3u l=0.1u
.ends OAI21X2

* Spice subcircuit definition for OAI21X4




.subckt OAI21X4 Y / A0 A1 B0
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n0 B0 Y VSS nmos1v w=1.72u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n1 A1 Y VDD pmos1v w=2.6u l=0.1u
mp2 Y B0 VDD VDD pmos1v w=2.6u l=0.1u
.ends OAI21X4

* Spice subcircuit definition for OAI21XL




.subckt OAI21XL Y / A0 A1 B0
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n0 B0 Y VSS nmos1v w=0.24u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1 Y VDD pmos1v w=0.36u l=0.1u
mp2 Y B0 VDD VDD pmos1v w=0.36u l=0.1u
.ends OAI21XL

* Spice subcircuit definition for OAI221X1




.subckt OAI221X1 Y / A0 A1 B0 B1 C0
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n0 B0 n1 VSS nmos1v w=0.43u l=0.1u
mn3 n0 B1 n1 VSS nmos1v w=0.43u l=0.1u
mn4 n1 C0 Y VSS nmos1v w=0.43u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n2 A1 Y VDD pmos1v w=0.65u l=0.1u
mp2 n3 B0 VDD VDD pmos1v w=0.65u l=0.1u
mp3 n3 B1 Y VDD pmos1v w=0.65u l=0.1u
mp4 Y C0 VDD VDD pmos1v w=0.65u l=0.1u
.ends OAI221X1

* Spice subcircuit definition for OAI221X2




.subckt OAI221X2 Y / A0 A1 B0 B1 C0
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.86u l=0.1u
mn2 n0 B0 n1 VSS nmos1v w=0.86u l=0.1u
mn3 n0 B1 n1 VSS nmos1v w=0.86u l=0.1u
mn4 n1 C0 Y VSS nmos1v w=0.86u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n2 A1 Y VDD pmos1v w=1.3u l=0.1u
mp2 n3 B0 VDD VDD pmos1v w=1.3u l=0.1u
mp3 n3 B1 Y VDD pmos1v w=1.3u l=0.1u
mp4 Y C0 VDD VDD pmos1v w=1.3u l=0.1u
.ends OAI221X2

* Spice subcircuit definition for OAI221X4




.subckt OAI221X4 Y / A0 A1 B0 B1 C0
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n0 B0 n1 VSS nmos1v w=1.72u l=0.1u
mn3 n0 B1 n1 VSS nmos1v w=1.72u l=0.1u
mn4 n1 C0 Y VSS nmos1v w=1.72u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n2 A1 Y VDD pmos1v w=2.6u l=0.1u
mp2 n3 B0 VDD VDD pmos1v w=2.6u l=0.1u
mp3 n3 B1 Y VDD pmos1v w=2.6u l=0.1u
mp4 Y C0 VDD VDD pmos1v w=2.6u l=0.1u
.ends OAI221X4

* Spice subcircuit definition for OAI221XL




.subckt OAI221XL Y / A0 A1 B0 B1 C0
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n0 B0 n1 VSS nmos1v w=0.24u l=0.1u
mn3 n0 B1 n1 VSS nmos1v w=0.24u l=0.1u
mn4 n1 C0 Y VSS nmos1v w=0.24u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 A1 Y VDD pmos1v w=0.36u l=0.1u
mp2 n3 B0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 B1 Y VDD pmos1v w=0.36u l=0.1u
mp4 Y C0 VDD VDD pmos1v w=0.36u l=0.1u
.ends OAI221XL

* Spice subcircuit definition for OAI222X1




.subckt OAI222X1 Y / A0 A1 B0 B1 C0 C1
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n0 B0 n1 VSS nmos1v w=0.43u l=0.1u
mn3 n0 B1 n1 VSS nmos1v w=0.43u l=0.1u
mn4 n1 C0 Y VSS nmos1v w=0.43u l=0.1u
mn5 n1 C1 Y VSS nmos1v w=0.43u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n2 A1 Y VDD pmos1v w=0.65u l=0.1u
mp2 n3 B0 VDD VDD pmos1v w=0.65u l=0.1u
mp3 n3 B1 Y VDD pmos1v w=0.65u l=0.1u
mp4 n4 C0 VDD VDD pmos1v w=0.65u l=0.1u
mp5 n4 C1 Y VDD pmos1v w=0.65u l=0.1u
.ends OAI222X1

* Spice subcircuit definition for OAI222X2




.subckt OAI222X2 Y / A0 A1 B0 B1 C0 C1
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.86u l=0.1u
mn2 n0 B0 n1 VSS nmos1v w=0.86u l=0.1u
mn3 n0 B1 n1 VSS nmos1v w=0.86u l=0.1u
mn4 n1 C0 Y VSS nmos1v w=0.86u l=0.1u
mn5 n1 C1 Y VSS nmos1v w=0.86u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n2 A1 Y VDD pmos1v w=1.3u l=0.1u
mp2 n3 B0 VDD VDD pmos1v w=1.3u l=0.1u
mp3 n3 B1 Y VDD pmos1v w=1.3u l=0.1u
mp4 n4 C0 VDD VDD pmos1v w=1.3u l=0.1u
mp5 n4 C1 Y VDD pmos1v w=1.3u l=0.1u
.ends OAI222X2

* Spice subcircuit definition for OAI222X4




.subckt OAI222X4 Y / A0 A1 B0 B1 C0 C1
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n0 B0 n1 VSS nmos1v w=1.72u l=0.1u
mn3 n0 B1 n1 VSS nmos1v w=1.72u l=0.1u
mn4 n1 C0 Y VSS nmos1v w=1.72u l=0.1u
mn5 n1 C1 Y VSS nmos1v w=1.72u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n2 A1 Y VDD pmos1v w=2.6u l=0.1u
mp2 n3 B0 VDD VDD pmos1v w=2.6u l=0.1u
mp3 n3 B1 Y VDD pmos1v w=2.6u l=0.1u
mp4 n4 C0 VDD VDD pmos1v w=2.6u l=0.1u
mp5 n4 C1 Y VDD pmos1v w=2.6u l=0.1u
.ends OAI222X4

* Spice subcircuit definition for OAI222XL




.subckt OAI222XL Y / A0 A1 B0 B1 C0 C1
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n0 B0 n1 VSS nmos1v w=0.24u l=0.1u
mn3 n0 B1 n1 VSS nmos1v w=0.24u l=0.1u
mn4 n1 C0 Y VSS nmos1v w=0.24u l=0.1u
mn5 n1 C1 Y VSS nmos1v w=0.24u l=0.1u
mp0 n2 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 A1 Y VDD pmos1v w=0.36u l=0.1u
mp2 n3 B0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 B1 Y VDD pmos1v w=0.36u l=0.1u
mp4 n4 C0 VDD VDD pmos1v w=0.36u l=0.1u
mp5 n4 C1 Y VDD pmos1v w=0.36u l=0.1u
.ends OAI222XL

* Spice subcircuit definition for OAI22X1




.subckt OAI22X1 Y / A0 A1 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n0 B0 Y VSS nmos1v w=0.43u l=0.1u
mn3 n0 B1 Y VSS nmos1v w=0.43u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 A1 Y VDD pmos1v w=0.65u l=0.1u
mp2 n2 B0 VDD VDD pmos1v w=0.65u l=0.1u
mp3 n2 B1 Y VDD pmos1v w=0.65u l=0.1u
.ends OAI22X1

* Spice subcircuit definition for OAI22X2




.subckt OAI22X2 Y / A0 A1 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.86u l=0.1u
mn2 n0 B0 Y VSS nmos1v w=0.86u l=0.1u
mn3 n0 B1 Y VSS nmos1v w=0.86u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n1 A1 Y VDD pmos1v w=1.3u l=0.1u
mp2 n2 B0 VDD VDD pmos1v w=1.3u l=0.1u
mp3 n2 B1 Y VDD pmos1v w=1.3u l=0.1u
.ends OAI22X2

* Spice subcircuit definition for OAI22X4




.subckt OAI22X4 Y / A0 A1 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n0 B0 Y VSS nmos1v w=1.72u l=0.1u
mn3 n0 B1 Y VSS nmos1v w=1.72u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n1 A1 Y VDD pmos1v w=2.6u l=0.1u
mp2 n2 B0 VDD VDD pmos1v w=2.6u l=0.1u
mp3 n2 B1 Y VDD pmos1v w=2.6u l=0.1u
.ends OAI22X4

* Spice subcircuit definition for OAI22XL




.subckt OAI22XL Y / A0 A1 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n0 B0 Y VSS nmos1v w=0.24u l=0.1u
mn3 n0 B1 Y VSS nmos1v w=0.24u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1 Y VDD pmos1v w=0.36u l=0.1u
mp2 n2 B0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n2 B1 Y VDD pmos1v w=0.36u l=0.1u
.ends OAI22XL

* Spice subcircuit definition for OAI2BB1X1




.subckt OAI2BB1X1 Y / A0N A1N B0
mn0 n1 A0N VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1N n0 VSS nmos1v w=0.24u l=0.1u
mn2 n2 B0 VSS VSS nmos1v w=0.43u l=0.1u
mn3 n2 n0 Y VSS nmos1v w=0.43u l=0.1u
mp0 n0 A0N VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 A1N VDD VDD pmos1v w=0.36u l=0.1u
mp2 Y B0 VDD VDD pmos1v w=0.65u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends OAI2BB1X1

* Spice subcircuit definition for OAI2BB1X2




.subckt OAI2BB1X2 Y / A0N A1N B0
mn0 n1 A0N VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1N n0 VSS nmos1v w=0.24u l=0.1u
mn2 n2 B0 VSS VSS nmos1v w=0.86u l=0.1u
mn3 n2 n0 Y VSS nmos1v w=0.86u l=0.1u
mp0 n0 A0N VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 A1N VDD VDD pmos1v w=0.36u l=0.1u
mp2 Y B0 VDD VDD pmos1v w=1.3u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends OAI2BB1X2

* Spice subcircuit definition for OAI2BB1X4




.subckt OAI2BB1X4 Y / A0N A1N B0
mn0 n1 A0N VSS VSS nmos1v w=0.43u l=0.1u
mn1 n1 A1N n0 VSS nmos1v w=0.43u l=0.1u
mn2 n2 B0 VSS VSS nmos1v w=1.72u l=0.1u
mn3 n2 n0 Y VSS nmos1v w=1.72u l=0.1u
mp0 n0 A0N VDD VDD pmos1v w=0.65u l=0.1u
mp1 n0 A1N VDD VDD pmos1v w=0.65u l=0.1u
mp2 Y B0 VDD VDD pmos1v w=2.6u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends OAI2BB1X4

* Spice subcircuit definition for OAI2BB1XL




.subckt OAI2BB1XL Y / A0N A1N B0
mn0 n1 A0N VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1N n0 VSS nmos1v w=0.24u l=0.1u
mn2 n2 B0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 n0 Y VSS nmos1v w=0.24u l=0.1u
mp0 n0 A0N VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 A1N VDD VDD pmos1v w=0.36u l=0.1u
mp2 Y B0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
.ends OAI2BB1XL

* Spice subcircuit definition for OAI2BB2X1




.subckt OAI2BB2X1 Y / A0N A1N B0 B1
mn0 n0 A0N VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1N VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=0.43u l=0.1u
mn3 n2 n1 VSS VSS nmos1v w=0.43u l=0.1u
mn4 n2 B0 Y VSS nmos1v w=0.43u l=0.1u
mn5 n2 B1 Y VSS nmos1v w=0.43u l=0.1u
mp0 n0 A0N VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1N VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 n0 VDD VDD pmos1v w=0.65u l=0.1u
mp3 n3 n1 Y VDD pmos1v w=0.65u l=0.1u
mp4 n4 B0 VDD VDD pmos1v w=0.65u l=0.1u
mp5 n4 B1 Y VDD pmos1v w=0.65u l=0.1u
.ends OAI2BB2X1

* Spice subcircuit definition for OAI2BB2X2




.subckt OAI2BB2X2 Y / A0N A1N B0 B1
mn0 n0 A0N VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1N VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=0.86u l=0.1u
mn3 n2 n1 VSS VSS nmos1v w=0.86u l=0.1u
mn4 n2 B0 Y VSS nmos1v w=0.86u l=0.1u
mn5 n2 B1 Y VSS nmos1v w=0.86u l=0.1u
mp0 n0 A0N VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1N VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 n0 VDD VDD pmos1v w=1.3u l=0.1u
mp3 n3 n1 Y VDD pmos1v w=1.3u l=0.1u
mp4 n4 B0 VDD VDD pmos1v w=1.3u l=0.1u
mp5 n4 B1 Y VDD pmos1v w=1.3u l=0.1u
.ends OAI2BB2X2

* Spice subcircuit definition for OAI2BB2X4




.subckt OAI2BB2X4 Y / A0N A1N B0 B1
mn0 n0 A0N VSS VSS nmos1v w=0.43u l=0.1u
mn1 n1 A1N VSS VSS nmos1v w=0.43u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=1.72u l=0.1u
mn3 n2 n1 VSS VSS nmos1v w=1.72u l=0.1u
mn4 n2 B0 Y VSS nmos1v w=1.72u l=0.1u
mn5 n2 B1 Y VSS nmos1v w=1.72u l=0.1u
mp0 n0 A0N VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 A1N VDD VDD pmos1v w=0.65u l=0.1u
mp2 n3 n0 VDD VDD pmos1v w=2.6u l=0.1u
mp3 n3 n1 Y VDD pmos1v w=2.6u l=0.1u
mp4 n4 B0 VDD VDD pmos1v w=2.6u l=0.1u
mp5 n4 B1 Y VDD pmos1v w=2.6u l=0.1u
.ends OAI2BB2X4

* Spice subcircuit definition for OAI2BB2XL




.subckt OAI2BB2XL Y / A0N A1N B0 B1
mn0 n0 A0N VSS VSS nmos1v w=0.24u l=0.1u
mn1 n1 A1N VSS VSS nmos1v w=0.24u l=0.1u
mn2 n2 n0 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n2 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn4 n2 B0 Y VSS nmos1v w=0.24u l=0.1u
mn5 n2 B1 Y VSS nmos1v w=0.24u l=0.1u
mp0 n0 A0N VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1N VDD VDD pmos1v w=0.36u l=0.1u
mp2 n3 n0 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n3 n1 Y VDD pmos1v w=0.36u l=0.1u
mp4 n4 B0 VDD VDD pmos1v w=0.36u l=0.1u
mp5 n4 B1 Y VDD pmos1v w=0.36u l=0.1u
.ends OAI2BB2XL

* Spice subcircuit definition for OAI31X1




.subckt OAI31X1 Y / A0 A1 A2 B0
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n0 A2 VSS VSS nmos1v w=0.43u l=0.1u
mn3 n0 B0 Y VSS nmos1v w=0.43u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 A1 n2 VDD pmos1v w=0.65u l=0.1u
mp2 n2 A2 Y VDD pmos1v w=0.65u l=0.1u
mp3 Y B0 VDD VDD pmos1v w=0.65u l=0.1u
.ends OAI31X1

* Spice subcircuit definition for OAI31X2




.subckt OAI31X2 Y / A0 A1 A2 B0
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.86u l=0.1u
mn2 n0 A2 VSS VSS nmos1v w=0.86u l=0.1u
mn3 n0 B0 Y VSS nmos1v w=0.86u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n1 A1 n2 VDD pmos1v w=1.3u l=0.1u
mp2 n2 A2 Y VDD pmos1v w=1.3u l=0.1u
mp3 Y B0 VDD VDD pmos1v w=1.3u l=0.1u
.ends OAI31X2

* Spice subcircuit definition for OAI31X4




.subckt OAI31X4 Y / A0 A1 A2 B0
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n0 A2 VSS VSS nmos1v w=1.72u l=0.1u
mn3 n0 B0 Y VSS nmos1v w=1.72u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n1 A1 n2 VDD pmos1v w=2.6u l=0.1u
mp2 n2 A2 Y VDD pmos1v w=2.6u l=0.1u
mp3 Y B0 VDD VDD pmos1v w=2.6u l=0.1u
.ends OAI31X4

* Spice subcircuit definition for OAI31XL




.subckt OAI31XL Y / A0 A1 A2 B0
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n0 A2 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n0 B0 Y VSS nmos1v w=0.24u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1 n2 VDD pmos1v w=0.36u l=0.1u
mp2 n2 A2 Y VDD pmos1v w=0.36u l=0.1u
mp3 Y B0 VDD VDD pmos1v w=0.36u l=0.1u
.ends OAI31XL

* Spice subcircuit definition for OAI32X1




.subckt OAI32X1 Y / A0 A1 A2 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n0 A2 VSS VSS nmos1v w=0.43u l=0.1u
mn3 n0 B0 Y VSS nmos1v w=0.43u l=0.1u
mn4 n0 B1 Y VSS nmos1v w=0.43u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 A1 n2 VDD pmos1v w=0.65u l=0.1u
mp2 n2 A2 Y VDD pmos1v w=0.65u l=0.1u
mp3 n3 B0 VDD VDD pmos1v w=0.65u l=0.1u
mp4 n3 B1 Y VDD pmos1v w=0.65u l=0.1u
.ends OAI32X1

* Spice subcircuit definition for OAI32X2




.subckt OAI32X2 Y / A0 A1 A2 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.86u l=0.1u
mn2 n0 A2 VSS VSS nmos1v w=0.86u l=0.1u
mn3 n0 B0 Y VSS nmos1v w=0.86u l=0.1u
mn4 n0 B1 Y VSS nmos1v w=0.86u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n1 A1 n2 VDD pmos1v w=1.3u l=0.1u
mp2 n2 A2 Y VDD pmos1v w=1.3u l=0.1u
mp3 n3 B0 VDD VDD pmos1v w=1.3u l=0.1u
mp4 n3 B1 Y VDD pmos1v w=1.3u l=0.1u
.ends OAI32X2

* Spice subcircuit definition for OAI32X4




.subckt OAI32X4 Y / A0 A1 A2 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n0 A2 VSS VSS nmos1v w=1.72u l=0.1u
mn3 n0 B0 Y VSS nmos1v w=1.72u l=0.1u
mn4 n0 B1 Y VSS nmos1v w=1.72u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n1 A1 n2 VDD pmos1v w=2.6u l=0.1u
mp2 n2 A2 Y VDD pmos1v w=2.6u l=0.1u
mp3 n3 B0 VDD VDD pmos1v w=2.6u l=0.1u
mp4 n3 B1 Y VDD pmos1v w=2.6u l=0.1u
.ends OAI32X4

* Spice subcircuit definition for OAI32XL




.subckt OAI32XL Y / A0 A1 A2 B0 B1
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n0 A2 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n0 B0 Y VSS nmos1v w=0.24u l=0.1u
mn4 n0 B1 Y VSS nmos1v w=0.24u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1 n2 VDD pmos1v w=0.36u l=0.1u
mp2 n2 A2 Y VDD pmos1v w=0.36u l=0.1u
mp3 n3 B0 VDD VDD pmos1v w=0.36u l=0.1u
mp4 n3 B1 Y VDD pmos1v w=0.36u l=0.1u
.ends OAI32XL

* Spice subcircuit definition for OAI33X1




.subckt OAI33X1 Y / A0 A1 A2 B0 B1 B2
mn0 n0 A0 VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.43u l=0.1u
mn2 n0 A2 VSS VSS nmos1v w=0.43u l=0.1u
mn3 n0 B0 Y VSS nmos1v w=0.43u l=0.1u
mn4 n0 B1 Y VSS nmos1v w=0.43u l=0.1u
mn5 n0 B2 Y VSS nmos1v w=0.43u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 A1 n2 VDD pmos1v w=0.65u l=0.1u
mp2 n2 A2 Y VDD pmos1v w=0.65u l=0.1u
mp3 n3 B0 VDD VDD pmos1v w=0.65u l=0.1u
mp4 n3 B1 n4 VDD pmos1v w=0.65u l=0.1u
mp5 n4 B2 Y VDD pmos1v w=0.65u l=0.1u
.ends OAI33X1

* Spice subcircuit definition for OAI33X2




.subckt OAI33X2 Y / A0 A1 A2 B0 B1 B2
mn0 n0 A0 VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.86u l=0.1u
mn2 n0 A2 VSS VSS nmos1v w=0.86u l=0.1u
mn3 n0 B0 Y VSS nmos1v w=0.86u l=0.1u
mn4 n0 B1 Y VSS nmos1v w=0.86u l=0.1u
mn5 n0 B2 Y VSS nmos1v w=0.86u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=1.3u l=0.1u
mp1 n1 A1 n2 VDD pmos1v w=1.3u l=0.1u
mp2 n2 A2 Y VDD pmos1v w=1.3u l=0.1u
mp3 n3 B0 VDD VDD pmos1v w=1.3u l=0.1u
mp4 n3 B1 n4 VDD pmos1v w=1.3u l=0.1u
mp5 n4 B2 Y VDD pmos1v w=1.3u l=0.1u
.ends OAI33X2

* Spice subcircuit definition for OAI33X4




.subckt OAI33X4 Y / A0 A1 A2 B0 B1 B2
mn0 n0 A0 VSS VSS nmos1v w=1.72u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=1.72u l=0.1u
mn2 n0 A2 VSS VSS nmos1v w=1.72u l=0.1u
mn3 n0 B0 Y VSS nmos1v w=1.72u l=0.1u
mn4 n0 B1 Y VSS nmos1v w=1.72u l=0.1u
mn5 n0 B2 Y VSS nmos1v w=1.72u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=2.6u l=0.1u
mp1 n1 A1 n2 VDD pmos1v w=2.6u l=0.1u
mp2 n2 A2 Y VDD pmos1v w=2.6u l=0.1u
mp3 n3 B0 VDD VDD pmos1v w=2.6u l=0.1u
mp4 n3 B1 n4 VDD pmos1v w=2.6u l=0.1u
mp5 n4 B2 Y VDD pmos1v w=2.6u l=0.1u
.ends OAI33X4

* Spice subcircuit definition for OAI33XL




.subckt OAI33XL Y / A0 A1 A2 B0 B1 B2
mn0 n0 A0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 A1 VSS VSS nmos1v w=0.24u l=0.1u
mn2 n0 A2 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n0 B0 Y VSS nmos1v w=0.24u l=0.1u
mn4 n0 B1 Y VSS nmos1v w=0.24u l=0.1u
mn5 n0 B2 Y VSS nmos1v w=0.24u l=0.1u
mp0 n1 A0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 A1 n2 VDD pmos1v w=0.36u l=0.1u
mp2 n2 A2 Y VDD pmos1v w=0.36u l=0.1u
mp3 n3 B0 VDD VDD pmos1v w=0.36u l=0.1u
mp4 n3 B1 n4 VDD pmos1v w=0.36u l=0.1u
mp5 n4 B2 Y VDD pmos1v w=0.36u l=0.1u
.ends OAI33XL

* Spice subcircuit definition for OR2X1




.subckt OR2X1 Y / A B
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B n0 VDD pmos1v w=0.36u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends OR2X1

* Spice subcircuit definition for OR2X2




.subckt OR2X2 Y / A B
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B n0 VDD pmos1v w=0.36u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends OR2X2

* Spice subcircuit definition for OR2X4




.subckt OR2X4 Y / A B
mn0 n0 A VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.43u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 B n0 VDD pmos1v w=0.65u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends OR2X4

* Spice subcircuit definition for OR2X6




.subckt OR2X6 Y / A B
mn0 n0 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.86u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=2.58u l=0.1u
mp0 n1 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n1 B n0 VDD pmos1v w=1.3u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=3.9u l=0.1u
.ends OR2X6

* Spice subcircuit definition for OR2X8




.subckt OR2X8 Y / A B
mn0 n0 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.86u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=3.44u l=0.1u
mp0 n1 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n1 B n0 VDD pmos1v w=1.3u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=5.2u l=0.1u
.ends OR2X8

* Spice subcircuit definition for OR2XL




.subckt OR2XL Y / A B
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B n0 VDD pmos1v w=0.36u l=0.1u
mp2 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
.ends OR2XL

* Spice subcircuit definition for OR3X1




.subckt OR3X1 Y / A B C
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n0 C VSS VSS nmos1v w=0.24u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B n2 VDD pmos1v w=0.36u l=0.1u
mp2 n2 C n0 VDD pmos1v w=0.36u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends OR3X1

* Spice subcircuit definition for OR3X2




.subckt OR3X2 Y / A B C
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n0 C VSS VSS nmos1v w=0.24u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B n2 VDD pmos1v w=0.36u l=0.1u
mp2 n2 C n0 VDD pmos1v w=0.36u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends OR3X2

* Spice subcircuit definition for OR3X4




.subckt OR3X4 Y / A B C
mn0 n0 A VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.43u l=0.1u
mn2 n0 C VSS VSS nmos1v w=0.43u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 B n2 VDD pmos1v w=0.65u l=0.1u
mp2 n2 C n0 VDD pmos1v w=0.65u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends OR3X4

* Spice subcircuit definition for OR3X6




.subckt OR3X6 Y / A B C
mn0 n0 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.86u l=0.1u
mn2 n0 C VSS VSS nmos1v w=0.86u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=2.58u l=0.1u
mp0 n1 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n1 B n2 VDD pmos1v w=1.3u l=0.1u
mp2 n2 C n0 VDD pmos1v w=1.3u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=3.9u l=0.1u
.ends OR3X6

* Spice subcircuit definition for OR3X8




.subckt OR3X8 Y / A B C
mn0 n0 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.86u l=0.1u
mn2 n0 C VSS VSS nmos1v w=0.86u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=3.44u l=0.1u
mp0 n1 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n1 B n2 VDD pmos1v w=1.3u l=0.1u
mp2 n2 C n0 VDD pmos1v w=1.3u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=5.2u l=0.1u
.ends OR3X8

* Spice subcircuit definition for OR3XL




.subckt OR3XL Y / A B C
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n0 C VSS VSS nmos1v w=0.24u l=0.1u
mn3 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B n2 VDD pmos1v w=0.36u l=0.1u
mp2 n2 C n0 VDD pmos1v w=0.36u l=0.1u
mp3 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
.ends OR3XL

* Spice subcircuit definition for OR4X1




.subckt OR4X1 Y / A B C D
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n0 C VSS VSS nmos1v w=0.24u l=0.1u
mn3 n0 D VSS VSS nmos1v w=0.24u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B n2 VDD pmos1v w=0.36u l=0.1u
mp2 n2 C n3 VDD pmos1v w=0.36u l=0.1u
mp3 n3 D n0 VDD pmos1v w=0.36u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends OR4X1

* Spice subcircuit definition for OR4X2




.subckt OR4X2 Y / A B C D
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n0 C VSS VSS nmos1v w=0.24u l=0.1u
mn3 n0 D VSS VSS nmos1v w=0.24u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B n2 VDD pmos1v w=0.36u l=0.1u
mp2 n2 C n3 VDD pmos1v w=0.36u l=0.1u
mp3 n3 D n0 VDD pmos1v w=0.36u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends OR4X2

* Spice subcircuit definition for OR4X4




.subckt OR4X4 Y / A B C D
mn0 n0 A VSS VSS nmos1v w=0.43u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.43u l=0.1u
mn2 n0 C VSS VSS nmos1v w=0.43u l=0.1u
mn3 n0 D VSS VSS nmos1v w=0.43u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.65u l=0.1u
mp1 n1 B n2 VDD pmos1v w=0.65u l=0.1u
mp2 n2 C n3 VDD pmos1v w=0.65u l=0.1u
mp3 n3 D n0 VDD pmos1v w=0.65u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends OR4X4

* Spice subcircuit definition for OR4X6




.subckt OR4X6 Y / A B C D
mn0 n0 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.86u l=0.1u
mn2 n0 C VSS VSS nmos1v w=0.86u l=0.1u
mn3 n0 D VSS VSS nmos1v w=0.86u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=2.58u l=0.1u
mp0 n1 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n1 B n2 VDD pmos1v w=1.3u l=0.1u
mp2 n2 C n3 VDD pmos1v w=1.3u l=0.1u
mp3 n3 D n0 VDD pmos1v w=1.3u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=3.9u l=0.1u
.ends OR4X6

* Spice subcircuit definition for OR4X8




.subckt OR4X8 Y / A B C D
mn0 n0 A VSS VSS nmos1v w=0.86u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.86u l=0.1u
mn2 n0 C VSS VSS nmos1v w=0.86u l=0.1u
mn3 n0 D VSS VSS nmos1v w=0.86u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=3.44u l=0.1u
mp0 n1 A VDD VDD pmos1v w=1.3u l=0.1u
mp1 n1 B n2 VDD pmos1v w=1.3u l=0.1u
mp2 n2 C n3 VDD pmos1v w=1.3u l=0.1u
mp3 n3 D n0 VDD pmos1v w=1.3u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=5.2u l=0.1u
.ends OR4X8

* Spice subcircuit definition for OR4XL




.subckt OR4XL Y / A B C D
mn0 n0 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n0 C VSS VSS nmos1v w=0.24u l=0.1u
mn3 n0 D VSS VSS nmos1v w=0.24u l=0.1u
mn4 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 B n2 VDD pmos1v w=0.36u l=0.1u
mp2 n2 C n3 VDD pmos1v w=0.36u l=0.1u
mp3 n3 D n0 VDD pmos1v w=0.36u l=0.1u
mp4 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
.ends OR4XL

* Spice subcircuit definition for SDFFHQX1




.subckt SDFFHQX1 Q / CK D SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
.ends SDFFHQX1

* Spice subcircuit definition for SDFFHQX2




.subckt SDFFHQX2 Q / CK D SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
.ends SDFFHQX2

* Spice subcircuit definition for SDFFHQX4




.subckt SDFFHQX4 Q / CK D SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
.ends SDFFHQX4

* Spice subcircuit definition for SDFFHQX8




.subckt SDFFHQX8 Q / CK D SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=1.29u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=3.44u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.95u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=5.2u l=0.1u
.ends SDFFHQX8

* Spice subcircuit definition for SDFFNSRX1




.subckt SDFFNSRX1 Q QN / CKN D RN SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKNb CKN VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKNbb CKNb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKNbb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKNb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKNb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKNbb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKNb CKN VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKNbb CKNb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKNb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKNbb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKNbb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKNb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
.ends SDFFNSRX1

* Spice subcircuit definition for SDFFNSRX2




.subckt SDFFNSRX2 Q QN / CKN D RN SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKNb CKN VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKNbb CKNb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKNbb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKNb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKNb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKNbb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKNb CKN VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKNbb CKNb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKNb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKNbb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKNbb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKNb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
.ends SDFFNSRX2

* Spice subcircuit definition for SDFFNSRX4




.subckt SDFFNSRX4 Q QN / CKN D RN SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKNb CKN VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKNbb CKNb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKNbb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKNb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKNb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKNbb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKNb CKN VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKNbb CKNb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKNb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKNbb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKNbb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKNb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
.ends SDFFNSRX4

* Spice subcircuit definition for SDFFNSRXL




.subckt SDFFNSRXL Q QN / CKN D RN SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKNb CKN VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKNbb CKNb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKNbb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKNb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKNb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKNbb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKNb CKN VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKNbb CKNb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKNb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKNbb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKNbb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKNb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
.ends SDFFNSRXL

* Spice subcircuit definition for SDFFQX1




.subckt SDFFQX1 Q / CK D SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
.ends SDFFQX1

* Spice subcircuit definition for SDFFQX2




.subckt SDFFQX2 Q / CK D SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
.ends SDFFQX2

* Spice subcircuit definition for SDFFQX4




.subckt SDFFQX4 Q / CK D SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
.ends SDFFQX4

* Spice subcircuit definition for SDFFQXL




.subckt SDFFQXL Q / CK D SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
.ends SDFFQXL

* Spice subcircuit definition for SDFFRHQX1




.subckt SDFFRHQX1 Q / CK D RN SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.34u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.34u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=0.34u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=0.34u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=0.52u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
.ends SDFFRHQX1

* Spice subcircuit definition for SDFFRHQX2




.subckt SDFFRHQX2 Q / CK D RN SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.34u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.34u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=0.34u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=0.34u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=0.52u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
.ends SDFFRHQX2

* Spice subcircuit definition for SDFFRHQX4




.subckt SDFFRHQX4 Q / CK D RN SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.34u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.34u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=0.68u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=0.68u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=1.04u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
.ends SDFFRHQX4

* Spice subcircuit definition for SDFFRHQX8




.subckt SDFFRHQX8 Q / CK D RN SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.34u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.34u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=1.29u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=1.29u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=3.44u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=1.95u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=1.95u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=5.2u l=0.1u
.ends SDFFRHQX8

* Spice subcircuit definition for SDFFRX1




.subckt SDFFRX1 Q QN / CK D RN SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.24u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.24u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=0.24u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=0.24u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=0.36u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
.ends SDFFRX1

* Spice subcircuit definition for SDFFRX2




.subckt SDFFRX2 Q QN / CK D RN SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.24u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.24u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=0.34u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=0.34u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=0.52u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
.ends SDFFRX2

* Spice subcircuit definition for SDFFRX4




.subckt SDFFRX4 Q QN / CK D RN SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.24u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.24u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=0.68u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=0.68u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=1.04u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
.ends SDFFRX4

* Spice subcircuit definition for SDFFRXL




.subckt SDFFRXL Q QN / CK D RN SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n27 RN VSS VSS nmos1v w=0.24u l=0.1u
mn36 n27 mout n25 VSS nmos1v w=0.24u l=0.1u
mn37 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 n35 RN VSS VSS nmos1v w=0.24u l=0.1u
mn46 n35 n30 qbint VSS nmos1v w=0.24u l=0.1u
mn50 n40 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n40 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 RN VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp37 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint RN VDD VDD pmos1v w=0.36u l=0.1u
mp46 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
.ends SDFFRXL

* Spice subcircuit definition for SDFFSHQX1




.subckt SDFFSHQX1 Q / CK D SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
.ends SDFFSHQX1

* Spice subcircuit definition for SDFFSHQX2




.subckt SDFFSHQX2 Q / CK D SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
.ends SDFFSHQX2

* Spice subcircuit definition for SDFFSHQX4




.subckt SDFFSHQX4 Q / CK D SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
.ends SDFFSHQX4

* Spice subcircuit definition for SDFFSHQX8




.subckt SDFFSHQX8 Q / CK D SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=1.29u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=3.44u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=1.95u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=5.2u l=0.1u
.ends SDFFSHQX8

* Spice subcircuit definition for SDFFSRHQX1




.subckt SDFFSRHQX1 Q / CK D RN SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.34u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.34u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.52u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
.ends SDFFSRHQX1

* Spice subcircuit definition for SDFFSRHQX2




.subckt SDFFSRHQX2 Q / CK D RN SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.34u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.34u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.52u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
.ends SDFFSRHQX2

* Spice subcircuit definition for SDFFSRHQX4




.subckt SDFFSRHQX4 Q / CK D RN SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.34u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.34u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.52u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
.ends SDFFSRHQX4

* Spice subcircuit definition for SDFFSRHQX8




.subckt SDFFSRHQX8 Q / CK D RN SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.43u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.43u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.43u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.34u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.34u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.34u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.34u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=1.29u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.34u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.34u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.34u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=3.44u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.65u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.65u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.65u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.52u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.52u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=1.95u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.52u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.52u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.52u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=5.2u l=0.1u
.ends SDFFSRHQX8

* Spice subcircuit definition for SDFFSRX1




.subckt SDFFSRX1 Q QN / CK D RN SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
.ends SDFFSRX1

* Spice subcircuit definition for SDFFSRX2




.subckt SDFFSRX2 Q QN / CK D RN SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
.ends SDFFSRX2

* Spice subcircuit definition for SDFFSRX4




.subckt SDFFSRX4 Q QN / CK D RN SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
.ends SDFFSRX4

* Spice subcircuit definition for SDFFSRXL




.subckt SDFFSRXL Q QN / CK D RN SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn22 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 RNb mout VSS nmos1v w=0.24u l=0.1u
mn32 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 RNb n40 VSS nmos1v w=0.24u l=0.1u
mn52 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn53 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp22 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 n26 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp32 n26 n20 mout VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n43 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp52 n43 qbint n41 VDD pmos1v w=0.36u l=0.1u
mp53 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
.ends SDFFSRXL

* Spice subcircuit definition for SDFFSX1




.subckt SDFFSX1 Q QN / CK D SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
.ends SDFFSX1

* Spice subcircuit definition for SDFFSX2




.subckt SDFFSX2 Q QN / CK D SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
.ends SDFFSX2

* Spice subcircuit definition for SDFFSX4




.subckt SDFFSX4 Q QN / CK D SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
.ends SDFFSX4

* Spice subcircuit definition for SDFFSXL




.subckt SDFFSXL Q QN / CK D SE SI SN
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 n25 SN VSS VSS nmos1v w=0.24u l=0.1u
mn31 n25 n20 mout VSS nmos1v w=0.24u l=0.1u
mn35 n30 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n30 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n35 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n35 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n42 SN VSS VSS nmos1v w=0.24u l=0.1u
mn51 n42 qbint n40 VSS nmos1v w=0.24u l=0.1u
mn52 n40 CKb n35 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout SN VDD VDD pmos1v w=0.36u l=0.1u
mp31 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n31 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n31 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n35 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n35 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n41 SN VDD VDD pmos1v w=0.36u l=0.1u
mp51 n41 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp52 n41 CKbb n35 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
.ends SDFFSXL

* Spice subcircuit definition for SDFFTRX1




.subckt SDFFTRX1 Q QN / CK D RN SE SI
mn0 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 D Db VSS nmos1v w=0.24u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 Db SEb Dbp VSS nmos1v w=0.24u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.24u l=0.1u
mn13 n10 SE Dbp VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dbp CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mp0 Db RN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 Db SE Dbp VDD pmos1v w=0.36u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.36u l=0.1u
mp13 n11 SEb Dbp VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dbp CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
.ends SDFFTRX1

* Spice subcircuit definition for SDFFTRX2




.subckt SDFFTRX2 Q QN / CK D RN SE SI
mn0 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 D Db VSS nmos1v w=0.24u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 Db SEb Dbp VSS nmos1v w=0.24u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.24u l=0.1u
mn13 n10 SE Dbp VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dbp CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mp0 Db RN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 Db SE Dbp VDD pmos1v w=0.36u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.36u l=0.1u
mp13 n11 SEb Dbp VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dbp CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
.ends SDFFTRX2

* Spice subcircuit definition for SDFFTRX4




.subckt SDFFTRX4 Q QN / CK D RN SE SI
mn0 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 D Db VSS nmos1v w=0.24u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 Db SEb Dbp VSS nmos1v w=0.24u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.24u l=0.1u
mn13 n10 SE Dbp VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dbp CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mp0 Db RN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 Db SE Dbp VDD pmos1v w=0.36u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.36u l=0.1u
mp13 n11 SEb Dbp VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dbp CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
.ends SDFFTRX4

* Spice subcircuit definition for SDFFTRXL




.subckt SDFFTRXL Q QN / CK D RN SE SI
mn0 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 D Db VSS nmos1v w=0.24u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 Db SEb Dbp VSS nmos1v w=0.24u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.24u l=0.1u
mn13 n10 SE Dbp VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dbp CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mp0 Db RN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 Db SE Dbp VDD pmos1v w=0.36u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.36u l=0.1u
mp13 n11 SEb Dbp VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dbp CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
.ends SDFFTRXL

* Spice subcircuit definition for SDFFX1




.subckt SDFFX1 Q QN / CK D SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
.ends SDFFX1

* Spice subcircuit definition for SDFFX2




.subckt SDFFX2 Q QN / CK D SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
.ends SDFFX2

* Spice subcircuit definition for SDFFX4




.subckt SDFFX4 Q QN / CK D SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
.ends SDFFX4

* Spice subcircuit definition for SDFFXL




.subckt SDFFXL Q QN / CK D SE SI
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 D VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Db VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Db CKb n20 VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 D VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Db VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Db CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
.ends SDFFXL

* Spice subcircuit definition for SEDFFHQX1




.subckt SEDFFHQX1 Q / CK D E SE SI
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 qint VSS VSS nmos1v w=0.43u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 Db SEb Dbp VSS nmos1v w=0.43u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.43u l=0.1u
mn13 n10 SE Dbp VSS nmos1v w=0.43u l=0.1u
mn2 n0 Eb Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dbp CKb n20 VSS nmos1v w=0.34u l=0.1u
mn3 n2 D VSS VSS nmos1v w=0.43u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn4 n2 E Db VSS nmos1v w=0.43u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.34u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 qint VDD VDD pmos1v w=0.65u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 Db SE Dbp VDD pmos1v w=0.65u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.65u l=0.1u
mp13 n11 SEb Dbp VDD pmos1v w=0.65u l=0.1u
mp2 n1 E Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dbp CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp3 n3 D VDD VDD pmos1v w=0.65u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp4 n3 Eb Db VDD pmos1v w=0.65u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.52u l=0.1u
.ends SEDFFHQX1

* Spice subcircuit definition for SEDFFHQX2




.subckt SEDFFHQX2 Q / CK D E SE SI
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 qint VSS VSS nmos1v w=0.43u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 Db SEb Dbp VSS nmos1v w=0.43u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.43u l=0.1u
mn13 n10 SE Dbp VSS nmos1v w=0.43u l=0.1u
mn2 n0 Eb Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dbp CKb n20 VSS nmos1v w=0.34u l=0.1u
mn3 n2 D VSS VSS nmos1v w=0.43u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn4 n2 E Db VSS nmos1v w=0.43u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.43u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.34u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 qint VDD VDD pmos1v w=0.65u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 Db SE Dbp VDD pmos1v w=0.65u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.65u l=0.1u
mp13 n11 SEb Dbp VDD pmos1v w=0.65u l=0.1u
mp2 n1 E Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dbp CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp3 n3 D VDD VDD pmos1v w=0.65u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp4 n3 Eb Db VDD pmos1v w=0.65u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.65u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.52u l=0.1u
.ends SEDFFHQX2

* Spice subcircuit definition for SEDFFHQX4




.subckt SEDFFHQX4 Q / CK D E SE SI
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 qint VSS VSS nmos1v w=0.43u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 Db SEb Dbp VSS nmos1v w=0.43u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.43u l=0.1u
mn13 n10 SE Dbp VSS nmos1v w=0.43u l=0.1u
mn2 n0 Eb Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dbp CKb n20 VSS nmos1v w=0.34u l=0.1u
mn3 n2 D VSS VSS nmos1v w=0.43u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn4 n2 E Db VSS nmos1v w=0.43u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 qint VDD VDD pmos1v w=0.65u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 Db SE Dbp VDD pmos1v w=0.65u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.65u l=0.1u
mp13 n11 SEb Dbp VDD pmos1v w=0.65u l=0.1u
mp2 n1 E Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dbp CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp3 n3 D VDD VDD pmos1v w=0.65u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp4 n3 Eb Db VDD pmos1v w=0.65u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
.ends SEDFFHQX4

* Spice subcircuit definition for SEDFFHQX8




.subckt SEDFFHQX8 Q / CK D E SE SI
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 qint VSS VSS nmos1v w=0.43u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 Db SEb Dbp VSS nmos1v w=0.43u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.43u l=0.1u
mn13 n10 SE Dbp VSS nmos1v w=0.43u l=0.1u
mn2 n0 Eb Db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dbp CKb n20 VSS nmos1v w=0.34u l=0.1u
mn3 n2 D VSS VSS nmos1v w=0.43u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn4 n2 E Db VSS nmos1v w=0.43u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=1.29u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=3.44u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.86u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 qint VDD VDD pmos1v w=0.65u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 Db SE Dbp VDD pmos1v w=0.65u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.65u l=0.1u
mp13 n11 SEb Dbp VDD pmos1v w=0.65u l=0.1u
mp2 n1 E Db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dbp CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp3 n3 D VDD VDD pmos1v w=0.65u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp4 n3 Eb Db VDD pmos1v w=0.65u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.95u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=5.2u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=1.3u l=0.1u
.ends SEDFFHQX8

* Spice subcircuit definition for SEDFFTRX1




.subckt SEDFFTRX1 Q QN / CK D E RN SE SI
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 Db D VSS VSS nmos1v w=0.24u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 Dp VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Dpb VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Dpb VSS nmos1v w=0.24u l=0.1u
mn2 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dpb CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 Dp RNb VSS VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn4 n0 Eb VSS VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn5 n0 qbint Dp VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mn6 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn7 n1 Db Dp VSS nmos1v w=0.24u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 Dp VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Dpb VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Dpb VDD pmos1v w=0.36u l=0.1u
mp2 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dpb CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n2 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp4 n2 Eb n3 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp5 n2 qbint n3 VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
mp6 n3 E Dp VDD pmos1v w=0.36u l=0.1u
mp7 n3 Db Dp VDD pmos1v w=0.36u l=0.1u
.ends SEDFFTRX1

* Spice subcircuit definition for SEDFFTRX2




.subckt SEDFFTRX2 Q QN / CK D E RN SE SI
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 Db D VSS VSS nmos1v w=0.24u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 Dp VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Dpb VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Dpb VSS nmos1v w=0.24u l=0.1u
mn2 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dpb CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 Dp RNb VSS VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn4 n0 Eb VSS VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn5 n0 qbint Dp VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mn6 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn7 n1 Db Dp VSS nmos1v w=0.24u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 Dp VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Dpb VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Dpb VDD pmos1v w=0.36u l=0.1u
mp2 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dpb CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n2 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp4 n2 Eb n3 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp5 n2 qbint n3 VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
mp6 n3 E Dp VDD pmos1v w=0.36u l=0.1u
mp7 n3 Db Dp VDD pmos1v w=0.36u l=0.1u
.ends SEDFFTRX2

* Spice subcircuit definition for SEDFFTRX4




.subckt SEDFFTRX4 Q QN / CK D E RN SE SI
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 Db D VSS VSS nmos1v w=0.24u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 Dp VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Dpb VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Dpb VSS nmos1v w=0.24u l=0.1u
mn2 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dpb CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 Dp RNb VSS VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn4 n0 Eb VSS VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn5 n0 qbint Dp VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mn6 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn7 n1 Db Dp VSS nmos1v w=0.24u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 Dp VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Dpb VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Dpb VDD pmos1v w=0.36u l=0.1u
mp2 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dpb CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n2 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp4 n2 Eb n3 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp5 n2 qbint n3 VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
mp6 n3 E Dp VDD pmos1v w=0.36u l=0.1u
mp7 n3 Db Dp VDD pmos1v w=0.36u l=0.1u
.ends SEDFFTRX4

* Spice subcircuit definition for SEDFFTRXL




.subckt SEDFFTRXL Q QN / CK D E RN SE SI
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 Db D VSS VSS nmos1v w=0.24u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 Dp VSS VSS nmos1v w=0.24u l=0.1u
mn12 n10 SEb Dpb VSS nmos1v w=0.24u l=0.1u
mn13 n12 SI VSS VSS nmos1v w=0.24u l=0.1u
mn14 n12 SE Dpb VSS nmos1v w=0.24u l=0.1u
mn2 RNb RN VSS VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dpb CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 Dp RNb VSS VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn4 n0 Eb VSS VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn5 n0 qbint Dp VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn7 n1 Db Dp VSS nmos1v w=0.24u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 Db D VDD VDD pmos1v w=0.36u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 n11 Dp VDD VDD pmos1v w=0.36u l=0.1u
mp12 n11 SE Dpb VDD pmos1v w=0.36u l=0.1u
mp13 n13 SI VDD VDD pmos1v w=0.36u l=0.1u
mp14 n13 SEb Dpb VDD pmos1v w=0.36u l=0.1u
mp2 RNb RN VDD VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dpb CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n2 RNb VDD VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp4 n2 Eb n3 VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp5 n2 qbint n3 VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
mp6 n3 E Dp VDD pmos1v w=0.36u l=0.1u
mp7 n3 Db Dp VDD pmos1v w=0.36u l=0.1u
.ends SEDFFTRXL

* Spice subcircuit definition for SEDFFX1




.subckt SEDFFX1 Q QN / CK D E SE SI
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 qint VSS VSS nmos1v w=0.24u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 Db SEb Dbp VSS nmos1v w=0.24u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.24u l=0.1u
mn13 n10 SE Dbp VSS nmos1v w=0.24u l=0.1u
mn2 n0 Eb Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dbp CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 n2 D VSS VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn4 n2 E Db VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.43u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 qint VDD VDD pmos1v w=0.36u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 Db SE Dbp VDD pmos1v w=0.36u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.36u l=0.1u
mp13 n11 SEb Dbp VDD pmos1v w=0.36u l=0.1u
mp2 n1 E Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dbp CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n3 D VDD VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp4 n3 Eb Db VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.65u l=0.1u
.ends SEDFFX1

* Spice subcircuit definition for SEDFFX2




.subckt SEDFFX2 Q QN / CK D E SE SI
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 qint VSS VSS nmos1v w=0.24u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 Db SEb Dbp VSS nmos1v w=0.24u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.24u l=0.1u
mn13 n10 SE Dbp VSS nmos1v w=0.24u l=0.1u
mn2 n0 Eb Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dbp CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 n2 D VSS VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn4 n2 E Db VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.86u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 qint VDD VDD pmos1v w=0.36u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 Db SE Dbp VDD pmos1v w=0.36u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.36u l=0.1u
mp13 n11 SEb Dbp VDD pmos1v w=0.36u l=0.1u
mp2 n1 E Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dbp CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n3 D VDD VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp4 n3 Eb Db VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=1.3u l=0.1u
.ends SEDFFX2

* Spice subcircuit definition for SEDFFX4




.subckt SEDFFX4 Q QN / CK D E SE SI
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 qint VSS VSS nmos1v w=0.24u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 Db SEb Dbp VSS nmos1v w=0.24u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.24u l=0.1u
mn13 n10 SE Dbp VSS nmos1v w=0.24u l=0.1u
mn2 n0 Eb Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dbp CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 n2 D VSS VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn4 n2 E Db VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.43u l=0.1u
mn57 QN qint VSS VSS nmos1v w=1.72u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 qint VDD VDD pmos1v w=0.36u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 Db SE Dbp VDD pmos1v w=0.36u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.36u l=0.1u
mp13 n11 SEb Dbp VDD pmos1v w=0.36u l=0.1u
mp2 n1 E Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dbp CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n3 D VDD VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp4 n3 Eb Db VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.65u l=0.1u
mp57 QN qint VDD VDD pmos1v w=2.6u l=0.1u
.ends SEDFFX4

* Spice subcircuit definition for SEDFFXL




.subckt SEDFFXL Q QN / CK D E SE SI
mn0 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 qint VSS VSS nmos1v w=0.24u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 Db SEb Dbp VSS nmos1v w=0.24u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.24u l=0.1u
mn13 n10 SE Dbp VSS nmos1v w=0.24u l=0.1u
mn2 n0 Eb Db VSS nmos1v w=0.24u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 Dbp CKb n20 VSS nmos1v w=0.24u l=0.1u
mn3 n2 D VSS VSS nmos1v w=0.24u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.24u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.24u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.24u l=0.1u
mn4 n2 E Db VSS nmos1v w=0.24u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.24u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.24u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.24u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.24u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.24u l=0.1u
mn56 qint qbint VSS VSS nmos1v w=0.24u l=0.1u
mn57 QN qint VSS VSS nmos1v w=0.24u l=0.1u
mp0 Eb E VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 qint VDD VDD pmos1v w=0.36u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 Db SE Dbp VDD pmos1v w=0.36u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.36u l=0.1u
mp13 n11 SEb Dbp VDD pmos1v w=0.36u l=0.1u
mp2 n1 E Db VDD pmos1v w=0.36u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 Dbp CKbb n20 VDD pmos1v w=0.36u l=0.1u
mp3 n3 D VDD VDD pmos1v w=0.36u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.36u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.36u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.36u l=0.1u
mp4 n3 Eb Db VDD pmos1v w=0.36u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.36u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.36u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.36u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.36u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.36u l=0.1u
mp56 qint qbint VDD VDD pmos1v w=0.36u l=0.1u
mp57 QN qint VDD VDD pmos1v w=0.36u l=0.1u
.ends SEDFFXL

* Spice subcircuit definition for SMDFFHQX1




.subckt SMDFFHQX1 Q / CK D0 D1 S0 SE SI
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 D0 VSS VSS nmos1v w=0.43u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 db SEb dbp VSS nmos1v w=0.43u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.43u l=0.1u
mn13 n10 SE dbp VSS nmos1v w=0.43u l=0.1u
mn2 n0 S0b db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 dbp CKb n20 VSS nmos1v w=0.34u l=0.1u
mn3 n2 D1 VSS VSS nmos1v w=0.43u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn4 n2 S0 db VSS nmos1v w=0.43u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.34u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.43u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 D0 VDD VDD pmos1v w=0.65u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 db SE dbp VDD pmos1v w=0.65u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.65u l=0.1u
mp13 n11 SEb dbp VDD pmos1v w=0.65u l=0.1u
mp2 n1 S0 db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 dbp CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp3 n3 D1 VDD VDD pmos1v w=0.65u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp4 n3 S0b db VDD pmos1v w=0.65u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.52u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=0.65u l=0.1u
.ends SMDFFHQX1

* Spice subcircuit definition for SMDFFHQX2




.subckt SMDFFHQX2 Q / CK D0 D1 S0 SE SI
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 D0 VSS VSS nmos1v w=0.43u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 db SEb dbp VSS nmos1v w=0.43u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.43u l=0.1u
mn13 n10 SE dbp VSS nmos1v w=0.43u l=0.1u
mn2 n0 S0b db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 dbp CKb n20 VSS nmos1v w=0.34u l=0.1u
mn3 n2 D1 VSS VSS nmos1v w=0.43u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn4 n2 S0 db VSS nmos1v w=0.43u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.43u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=0.86u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 D0 VDD VDD pmos1v w=0.65u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 db SE dbp VDD pmos1v w=0.65u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.65u l=0.1u
mp13 n11 SEb dbp VDD pmos1v w=0.65u l=0.1u
mp2 n1 S0 db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 dbp CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp3 n3 D1 VDD VDD pmos1v w=0.65u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp4 n3 S0b db VDD pmos1v w=0.65u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=0.65u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=1.3u l=0.1u
.ends SMDFFHQX2

* Spice subcircuit definition for SMDFFHQX4




.subckt SMDFFHQX4 Q / CK D0 D1 S0 SE SI
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 D0 VSS VSS nmos1v w=0.43u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 db SEb dbp VSS nmos1v w=0.43u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.43u l=0.1u
mn13 n10 SE dbp VSS nmos1v w=0.43u l=0.1u
mn2 n0 S0b db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 dbp CKb n20 VSS nmos1v w=0.34u l=0.1u
mn3 n2 D1 VSS VSS nmos1v w=0.43u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn4 n2 S0 db VSS nmos1v w=0.43u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=0.68u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=1.72u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 D0 VDD VDD pmos1v w=0.65u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 db SE dbp VDD pmos1v w=0.65u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.65u l=0.1u
mp13 n11 SEb dbp VDD pmos1v w=0.65u l=0.1u
mp2 n1 S0 db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 dbp CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp3 n3 D1 VDD VDD pmos1v w=0.65u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp4 n3 S0b db VDD pmos1v w=0.65u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.04u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=2.6u l=0.1u
.ends SMDFFHQX4

* Spice subcircuit definition for SMDFFHQX8




.subckt SMDFFHQX8 Q / CK D0 D1 S0 SE SI
mn0 S0b S0 VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 D0 VSS VSS nmos1v w=0.43u l=0.1u
mn10 SEb SE VSS VSS nmos1v w=0.24u l=0.1u
mn11 db SEb dbp VSS nmos1v w=0.43u l=0.1u
mn12 n10 SI VSS VSS nmos1v w=0.43u l=0.1u
mn13 n10 SE dbp VSS nmos1v w=0.43u l=0.1u
mn2 n0 S0b db VSS nmos1v w=0.43u l=0.1u
mn20 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn21 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn25 dbp CKb n20 VSS nmos1v w=0.34u l=0.1u
mn3 n2 D1 VSS VSS nmos1v w=0.43u l=0.1u
mn30 mout n20 VSS VSS nmos1v w=0.34u l=0.1u
mn35 n25 mout VSS VSS nmos1v w=0.34u l=0.1u
mn36 n25 CKbb n20 VSS nmos1v w=0.34u l=0.1u
mn4 n2 S0 db VSS nmos1v w=0.43u l=0.1u
mn40 mout CKbb n30 VSS nmos1v w=0.34u l=0.1u
mn45 qbint n30 VSS VSS nmos1v w=1.29u l=0.1u
mn50 n35 qbint VSS VSS nmos1v w=0.34u l=0.1u
mn51 n35 CKb n30 VSS nmos1v w=0.34u l=0.1u
mn55 Q qbint VSS VSS nmos1v w=3.44u l=0.1u
mp0 S0b S0 VDD VDD pmos1v w=0.36u l=0.1u
mp1 n1 D0 VDD VDD pmos1v w=0.65u l=0.1u
mp10 SEb SE VDD VDD pmos1v w=0.36u l=0.1u
mp11 db SE dbp VDD pmos1v w=0.65u l=0.1u
mp12 n11 SI VDD VDD pmos1v w=0.65u l=0.1u
mp13 n11 SEb dbp VDD pmos1v w=0.65u l=0.1u
mp2 n1 S0 db VDD pmos1v w=0.65u l=0.1u
mp20 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp21 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp25 dbp CKbb n20 VDD pmos1v w=0.52u l=0.1u
mp3 n3 D1 VDD VDD pmos1v w=0.65u l=0.1u
mp30 mout n20 VDD VDD pmos1v w=0.52u l=0.1u
mp35 n26 mout VDD VDD pmos1v w=0.52u l=0.1u
mp36 n26 CKb n20 VDD pmos1v w=0.52u l=0.1u
mp4 n3 S0b db VDD pmos1v w=0.65u l=0.1u
mp40 mout CKb n30 VDD pmos1v w=0.52u l=0.1u
mp45 qbint n30 VDD VDD pmos1v w=1.95u l=0.1u
mp50 n36 qbint VDD VDD pmos1v w=0.52u l=0.1u
mp51 n36 CKbb n30 VDD pmos1v w=0.52u l=0.1u
mp55 Q qbint VDD VDD pmos1v w=5.2u l=0.1u
.ends SMDFFHQX8

* Spice subcircuit definition for TBUFX1




.subckt TBUFX1 Y / A OE
mn0 OEb OE VSS VSS nmos1v w=0.24u l=0.1u
mn1 non A VSS VSS nmos1v w=0.24u l=0.1u
mn2 non OEb VSS VSS nmos1v w=0.24u l=0.1u
mn3 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn4 n1 OE pon VSS nmos1v w=0.24u l=0.1u
mn5 Y non VSS VSS nmos1v w=0.43u l=0.1u
mp0 OEb OE VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp2 n0 OEb non VDD pmos1v w=0.36u l=0.1u
mp3 pon A VDD VDD pmos1v w=0.36u l=0.1u
mp4 pon OE VDD VDD pmos1v w=0.36u l=0.1u
mp5 Y pon VDD VDD pmos1v w=0.65u l=0.1u
.ends TBUFX1

* Spice subcircuit definition for TBUFX12




.subckt TBUFX12 Y / A OE
mn0 OEb OE VSS VSS nmos1v w=0.43u l=0.1u
mn1 non A VSS VSS nmos1v w=1.29u l=0.1u
mn2 non OEb VSS VSS nmos1v w=1.29u l=0.1u
mn3 n1 A VSS VSS nmos1v w=1.29u l=0.1u
mn4 n1 OE pon VSS nmos1v w=1.29u l=0.1u
mn5 Y non VSS VSS nmos1v w=5.16u l=0.1u
mp0 OEb OE VDD VDD pmos1v w=0.65u l=0.1u
mp1 n0 A VDD VDD pmos1v w=1.95u l=0.1u
mp2 n0 OEb non VDD pmos1v w=1.95u l=0.1u
mp3 pon A VDD VDD pmos1v w=1.95u l=0.1u
mp4 pon OE VDD VDD pmos1v w=1.95u l=0.1u
mp5 Y pon VDD VDD pmos1v w=7.8u l=0.1u
.ends TBUFX12

* Spice subcircuit definition for TBUFX16




.subckt TBUFX16 Y / A OE
mn0 OEb OE VSS VSS nmos1v w=0.43u l=0.1u
mn1 non A VSS VSS nmos1v w=1.72u l=0.1u
mn2 non OEb VSS VSS nmos1v w=1.72u l=0.1u
mn3 n1 A VSS VSS nmos1v w=1.72u l=0.1u
mn4 n1 OE pon VSS nmos1v w=1.72u l=0.1u
mn5 Y non VSS VSS nmos1v w=6.88u l=0.1u
mp0 OEb OE VDD VDD pmos1v w=0.65u l=0.1u
mp1 n0 A VDD VDD pmos1v w=2.6u l=0.1u
mp2 n0 OEb non VDD pmos1v w=2.6u l=0.1u
mp3 pon A VDD VDD pmos1v w=2.6u l=0.1u
mp4 pon OE VDD VDD pmos1v w=2.6u l=0.1u
mp5 Y pon VDD VDD pmos1v w=10.4u l=0.1u
.ends TBUFX16

* Spice subcircuit definition for TBUFX2




.subckt TBUFX2 Y / A OE
mn0 OEb OE VSS VSS nmos1v w=0.24u l=0.1u
mn1 non A VSS VSS nmos1v w=0.24u l=0.1u
mn2 non OEb VSS VSS nmos1v w=0.24u l=0.1u
mn3 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn4 n1 OE pon VSS nmos1v w=0.24u l=0.1u
mn5 Y non VSS VSS nmos1v w=0.86u l=0.1u
mp0 OEb OE VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp2 n0 OEb non VDD pmos1v w=0.36u l=0.1u
mp3 pon A VDD VDD pmos1v w=0.36u l=0.1u
mp4 pon OE VDD VDD pmos1v w=0.36u l=0.1u
mp5 Y pon VDD VDD pmos1v w=1.3u l=0.1u
.ends TBUFX2

* Spice subcircuit definition for TBUFX20




.subckt TBUFX20 Y / A OE
mn0 OEb OE VSS VSS nmos1v w=0.86u l=0.1u
mn1 non A VSS VSS nmos1v w=2.15u l=0.1u
mn2 non OEb VSS VSS nmos1v w=2.15u l=0.1u
mn3 n1 A VSS VSS nmos1v w=2.15u l=0.1u
mn4 n1 OE pon VSS nmos1v w=2.15u l=0.1u
mn5 Y non VSS VSS nmos1v w=8.6u l=0.1u
mp0 OEb OE VDD VDD pmos1v w=1.3u l=0.1u
mp1 n0 A VDD VDD pmos1v w=3.25u l=0.1u
mp2 n0 OEb non VDD pmos1v w=3.25u l=0.1u
mp3 pon A VDD VDD pmos1v w=3.25u l=0.1u
mp4 pon OE VDD VDD pmos1v w=3.25u l=0.1u
mp5 Y pon VDD VDD pmos1v w=13.0u l=0.1u
.ends TBUFX20

* Spice subcircuit definition for TBUFX3




.subckt TBUFX3 Y / A OE
mn0 OEb OE VSS VSS nmos1v w=0.24u l=0.1u
mn1 non A VSS VSS nmos1v w=0.43u l=0.1u
mn2 non OEb VSS VSS nmos1v w=0.43u l=0.1u
mn3 n1 A VSS VSS nmos1v w=0.43u l=0.1u
mn4 n1 OE pon VSS nmos1v w=0.43u l=0.1u
mn5 Y non VSS VSS nmos1v w=1.29u l=0.1u
mp0 OEb OE VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 A VDD VDD pmos1v w=0.65u l=0.1u
mp2 n0 OEb non VDD pmos1v w=0.65u l=0.1u
mp3 pon A VDD VDD pmos1v w=0.65u l=0.1u
mp4 pon OE VDD VDD pmos1v w=0.65u l=0.1u
mp5 Y pon VDD VDD pmos1v w=1.95u l=0.1u
.ends TBUFX3

* Spice subcircuit definition for TBUFX4




.subckt TBUFX4 Y / A OE
mn0 OEb OE VSS VSS nmos1v w=0.24u l=0.1u
mn1 non A VSS VSS nmos1v w=0.43u l=0.1u
mn2 non OEb VSS VSS nmos1v w=0.43u l=0.1u
mn3 n1 A VSS VSS nmos1v w=0.43u l=0.1u
mn4 n1 OE pon VSS nmos1v w=0.43u l=0.1u
mn5 Y non VSS VSS nmos1v w=1.72u l=0.1u
mp0 OEb OE VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 A VDD VDD pmos1v w=0.65u l=0.1u
mp2 n0 OEb non VDD pmos1v w=0.65u l=0.1u
mp3 pon A VDD VDD pmos1v w=0.65u l=0.1u
mp4 pon OE VDD VDD pmos1v w=0.65u l=0.1u
mp5 Y pon VDD VDD pmos1v w=2.6u l=0.1u
.ends TBUFX4

* Spice subcircuit definition for TBUFX6




.subckt TBUFX6 Y / A OE
mn0 OEb OE VSS VSS nmos1v w=0.24u l=0.1u
mn1 non A VSS VSS nmos1v w=0.86u l=0.1u
mn2 non OEb VSS VSS nmos1v w=0.86u l=0.1u
mn3 n1 A VSS VSS nmos1v w=0.86u l=0.1u
mn4 n1 OE pon VSS nmos1v w=0.86u l=0.1u
mn5 Y non VSS VSS nmos1v w=2.58u l=0.1u
mp0 OEb OE VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp2 n0 OEb non VDD pmos1v w=1.3u l=0.1u
mp3 pon A VDD VDD pmos1v w=1.3u l=0.1u
mp4 pon OE VDD VDD pmos1v w=1.3u l=0.1u
mp5 Y pon VDD VDD pmos1v w=3.9u l=0.1u
.ends TBUFX6

* Spice subcircuit definition for TBUFX8




.subckt TBUFX8 Y / A OE
mn0 OEb OE VSS VSS nmos1v w=0.24u l=0.1u
mn1 non A VSS VSS nmos1v w=0.86u l=0.1u
mn2 non OEb VSS VSS nmos1v w=0.86u l=0.1u
mn3 n1 A VSS VSS nmos1v w=0.86u l=0.1u
mn4 n1 OE pon VSS nmos1v w=0.86u l=0.1u
mn5 Y non VSS VSS nmos1v w=3.44u l=0.1u
mp0 OEb OE VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 A VDD VDD pmos1v w=1.3u l=0.1u
mp2 n0 OEb non VDD pmos1v w=1.3u l=0.1u
mp3 pon A VDD VDD pmos1v w=1.3u l=0.1u
mp4 pon OE VDD VDD pmos1v w=1.3u l=0.1u
mp5 Y pon VDD VDD pmos1v w=5.2u l=0.1u
.ends TBUFX8

* Spice subcircuit definition for TBUFXL




.subckt TBUFXL Y / A OE
mn0 OEb OE VSS VSS nmos1v w=0.24u l=0.1u
mn1 non A VSS VSS nmos1v w=0.24u l=0.1u
mn2 non OEb VSS VSS nmos1v w=0.24u l=0.1u
mn3 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn4 n1 OE pon VSS nmos1v w=0.24u l=0.1u
mn5 Y non VSS VSS nmos1v w=0.24u l=0.1u
mp0 OEb OE VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 A VDD VDD pmos1v w=0.36u l=0.1u
mp2 n0 OEb non VDD pmos1v w=0.36u l=0.1u
mp3 pon A VDD VDD pmos1v w=0.36u l=0.1u
mp4 pon OE VDD VDD pmos1v w=0.36u l=0.1u
mp5 Y pon VDD VDD pmos1v w=0.36u l=0.1u
.ends TBUFXL

* Spice subcircuit definition for TIEHI




.subckt TIEHI Y /
mn0 n0 n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends TIEHI

* Spice subcircuit definition for TIELO




.subckt TIELO Y /
mn0 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n0 n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends TIELO

* Spice subcircuit definition for TLATNCAX12




.subckt TLATNCAX12 ECK / CK E
mn0 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn1 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n0 VSS VSS nmos1v w=0.43u l=0.1u
mn15 n5 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 CKbb n0 VSS nmos1v w=0.24u l=0.1u
mn20 n10 Eint VSS VSS nmos1v w=1.29u l=0.1u
mn21 n10 CKbb ECKb VSS nmos1v w=1.29u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=5.16u l=0.1u
mn5 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 CKb n0 VSS nmos1v w=0.24u l=0.1u
mp0 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp1 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Eint n0 VDD VDD pmos1v w=0.65u l=0.1u
mp15 n6 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 CKb n0 VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=1.95u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=1.95u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=7.8u l=0.1u
mp5 n2 E VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 CKbb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATNCAX12

* Spice subcircuit definition for TLATNCAX16




.subckt TLATNCAX16 ECK / CK E
mn0 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn1 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n0 VSS VSS nmos1v w=0.68u l=0.1u
mn15 n5 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 CKbb n0 VSS nmos1v w=0.24u l=0.1u
mn20 n10 Eint VSS VSS nmos1v w=1.72u l=0.1u
mn21 n10 CKbb ECKb VSS nmos1v w=1.72u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=6.88u l=0.1u
mn5 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 CKb n0 VSS nmos1v w=0.24u l=0.1u
mp0 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp1 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Eint n0 VDD VDD pmos1v w=1.04u l=0.1u
mp15 n6 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 CKb n0 VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=2.6u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=2.6u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=10.4u l=0.1u
mp5 n2 E VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 CKbb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATNCAX16

* Spice subcircuit definition for TLATNCAX2




.subckt TLATNCAX2 ECK / CK E
mn0 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn1 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n0 VSS VSS nmos1v w=0.24u l=0.1u
mn15 n5 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 CKbb n0 VSS nmos1v w=0.24u l=0.1u
mn20 n10 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn21 n10 CKbb ECKb VSS nmos1v w=0.24u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=0.86u l=0.1u
mn5 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 CKb n0 VSS nmos1v w=0.24u l=0.1u
mp0 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp1 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Eint n0 VDD VDD pmos1v w=0.36u l=0.1u
mp15 n6 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 CKb n0 VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=0.36u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=0.36u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=1.3u l=0.1u
mp5 n2 E VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 CKbb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATNCAX2

* Spice subcircuit definition for TLATNCAX20




.subckt TLATNCAX20 ECK / CK E
mn0 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn1 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n0 VSS VSS nmos1v w=0.86u l=0.1u
mn15 n5 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 CKbb n0 VSS nmos1v w=0.24u l=0.1u
mn20 n10 Eint VSS VSS nmos1v w=2.15u l=0.1u
mn21 n10 CKbb ECKb VSS nmos1v w=2.15u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=8.6u l=0.1u
mn5 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 CKb n0 VSS nmos1v w=0.24u l=0.1u
mp0 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp1 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Eint n0 VDD VDD pmos1v w=1.3u l=0.1u
mp15 n6 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 CKb n0 VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=3.25u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=3.25u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=13.0u l=0.1u
mp5 n2 E VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 CKbb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATNCAX20

* Spice subcircuit definition for TLATNCAX3




.subckt TLATNCAX3 ECK / CK E
mn0 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn1 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n0 VSS VSS nmos1v w=0.24u l=0.1u
mn15 n5 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 CKbb n0 VSS nmos1v w=0.24u l=0.1u
mn20 n10 Eint VSS VSS nmos1v w=0.43u l=0.1u
mn21 n10 CKbb ECKb VSS nmos1v w=0.43u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=1.29u l=0.1u
mn5 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 CKb n0 VSS nmos1v w=0.24u l=0.1u
mp0 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp1 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Eint n0 VDD VDD pmos1v w=0.36u l=0.1u
mp15 n6 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 CKb n0 VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=0.65u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=0.65u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=1.95u l=0.1u
mp5 n2 E VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 CKbb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATNCAX3

* Spice subcircuit definition for TLATNCAX4




.subckt TLATNCAX4 ECK / CK E
mn0 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn1 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n0 VSS VSS nmos1v w=0.24u l=0.1u
mn15 n5 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 CKbb n0 VSS nmos1v w=0.24u l=0.1u
mn20 n10 Eint VSS VSS nmos1v w=0.43u l=0.1u
mn21 n10 CKbb ECKb VSS nmos1v w=0.43u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=1.72u l=0.1u
mn5 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 CKb n0 VSS nmos1v w=0.24u l=0.1u
mp0 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp1 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Eint n0 VDD VDD pmos1v w=0.36u l=0.1u
mp15 n6 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 CKb n0 VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=0.65u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=0.65u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=2.6u l=0.1u
mp5 n2 E VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 CKbb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATNCAX4

* Spice subcircuit definition for TLATNCAX6




.subckt TLATNCAX6 ECK / CK E
mn0 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn1 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n0 VSS VSS nmos1v w=0.34u l=0.1u
mn15 n5 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 CKbb n0 VSS nmos1v w=0.24u l=0.1u
mn20 n10 Eint VSS VSS nmos1v w=0.86u l=0.1u
mn21 n10 CKbb ECKb VSS nmos1v w=0.86u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=2.58u l=0.1u
mn5 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 CKb n0 VSS nmos1v w=0.24u l=0.1u
mp0 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp1 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Eint n0 VDD VDD pmos1v w=0.52u l=0.1u
mp15 n6 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 CKb n0 VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=1.3u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=1.3u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=3.9u l=0.1u
mp5 n2 E VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 CKbb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATNCAX6

* Spice subcircuit definition for TLATNCAX8




.subckt TLATNCAX8 ECK / CK E
mn0 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn1 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n0 VSS VSS nmos1v w=0.34u l=0.1u
mn15 n5 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 CKbb n0 VSS nmos1v w=0.24u l=0.1u
mn20 n10 Eint VSS VSS nmos1v w=0.86u l=0.1u
mn21 n10 CKbb ECKb VSS nmos1v w=0.86u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=3.44u l=0.1u
mn5 n1 E VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 CKb n0 VSS nmos1v w=0.24u l=0.1u
mp0 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp1 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Eint n0 VDD VDD pmos1v w=0.52u l=0.1u
mp15 n6 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 CKb n0 VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=1.3u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=1.3u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=5.2u l=0.1u
mp5 n2 E VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 CKbb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATNCAX8

* Spice subcircuit definition for TLATNSRX1




.subckt TLATNSRX1 Q QN / D GN RN SN
mn0 GNbp GN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn10 n10 SN VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 n5 Qint VSS nmos1v w=0.24u l=0.1u
mn15 n17 RN VSS VSS nmos1v w=0.24u l=0.1u
mn16 n17 Qint n15 VSS nmos1v w=0.24u l=0.1u
mn17 n15 GNbb n5 VSS nmos1v w=0.24u l=0.1u
mn2 n0 GNbp GNbb VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=0.43u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=0.43u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=0.43u l=0.1u
mn3 GNb GNbb VSS VSS nmos1v w=0.24u l=0.1u
mn5 n6 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n6 GNb n5 VSS nmos1v w=0.24u l=0.1u
mp0 GNbp GN VDD VDD pmos1v w=0.36u l=0.1u
mp1 GNbb RN VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint SN VDD VDD pmos1v w=0.36u l=0.1u
mp11 Qint n5 VDD VDD pmos1v w=0.36u l=0.1u
mp15 n16 RN VDD VDD pmos1v w=0.36u l=0.1u
mp16 n16 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp17 n16 GNb n5 VDD pmos1v w=0.36u l=0.1u
mp2 GNbb GNbp VDD VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=0.65u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=0.65u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=0.65u l=0.1u
mp3 GNb GNbb VDD VDD pmos1v w=0.36u l=0.1u
mp5 n7 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n7 GNbb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATNSRX1

* Spice subcircuit definition for TLATNSRX2




.subckt TLATNSRX2 Q QN / D GN RN SN
mn0 GNbp GN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn10 n10 SN VSS VSS nmos1v w=0.34u l=0.1u
mn11 n10 n5 Qint VSS nmos1v w=0.34u l=0.1u
mn15 n17 RN VSS VSS nmos1v w=0.24u l=0.1u
mn16 n17 Qint n15 VSS nmos1v w=0.24u l=0.1u
mn17 n15 GNbb n5 VSS nmos1v w=0.24u l=0.1u
mn2 n0 GNbp GNbb VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=0.86u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=0.86u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=0.86u l=0.1u
mn3 GNb GNbb VSS VSS nmos1v w=0.24u l=0.1u
mn5 n6 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n6 GNb n5 VSS nmos1v w=0.24u l=0.1u
mp0 GNbp GN VDD VDD pmos1v w=0.36u l=0.1u
mp1 GNbb RN VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint SN VDD VDD pmos1v w=0.52u l=0.1u
mp11 Qint n5 VDD VDD pmos1v w=0.52u l=0.1u
mp15 n16 RN VDD VDD pmos1v w=0.36u l=0.1u
mp16 n16 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp17 n16 GNb n5 VDD pmos1v w=0.36u l=0.1u
mp2 GNbb GNbp VDD VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=1.3u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=1.3u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=1.3u l=0.1u
mp3 GNb GNbb VDD VDD pmos1v w=0.36u l=0.1u
mp5 n7 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n7 GNbb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATNSRX2

* Spice subcircuit definition for TLATNSRX4




.subckt TLATNSRX4 Q QN / D GN RN SN
mn0 GNbp GN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn10 n10 SN VSS VSS nmos1v w=0.68u l=0.1u
mn11 n10 n5 Qint VSS nmos1v w=0.68u l=0.1u
mn15 n17 RN VSS VSS nmos1v w=0.24u l=0.1u
mn16 n17 Qint n15 VSS nmos1v w=0.24u l=0.1u
mn17 n15 GNbb n5 VSS nmos1v w=0.24u l=0.1u
mn2 n0 GNbp GNbb VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=1.72u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=1.72u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=1.72u l=0.1u
mn3 GNb GNbb VSS VSS nmos1v w=0.24u l=0.1u
mn5 n6 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n6 GNb n5 VSS nmos1v w=0.24u l=0.1u
mp0 GNbp GN VDD VDD pmos1v w=0.36u l=0.1u
mp1 GNbb RN VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint SN VDD VDD pmos1v w=1.04u l=0.1u
mp11 Qint n5 VDD VDD pmos1v w=1.04u l=0.1u
mp15 n16 RN VDD VDD pmos1v w=0.36u l=0.1u
mp16 n16 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp17 n16 GNb n5 VDD pmos1v w=0.36u l=0.1u
mp2 GNbb GNbp VDD VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=2.6u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=2.6u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=2.6u l=0.1u
mp3 GNb GNbb VDD VDD pmos1v w=0.36u l=0.1u
mp5 n7 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n7 GNbb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATNSRX4

* Spice subcircuit definition for TLATNSRXL




.subckt TLATNSRXL Q QN / D GN RN SN
mn0 GNbp GN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn10 n10 SN VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 n5 Qint VSS nmos1v w=0.24u l=0.1u
mn15 n17 RN VSS VSS nmos1v w=0.24u l=0.1u
mn16 n17 Qint n15 VSS nmos1v w=0.24u l=0.1u
mn17 n15 GNbb n5 VSS nmos1v w=0.24u l=0.1u
mn2 n0 GNbp GNbb VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=0.24u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=0.24u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=0.24u l=0.1u
mn3 GNb GNbb VSS VSS nmos1v w=0.24u l=0.1u
mn5 n6 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n6 GNb n5 VSS nmos1v w=0.24u l=0.1u
mp0 GNbp GN VDD VDD pmos1v w=0.36u l=0.1u
mp1 GNbb RN VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint SN VDD VDD pmos1v w=0.36u l=0.1u
mp11 Qint n5 VDD VDD pmos1v w=0.36u l=0.1u
mp15 n16 RN VDD VDD pmos1v w=0.36u l=0.1u
mp16 n16 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp17 n16 GNb n5 VDD pmos1v w=0.36u l=0.1u
mp2 GNbb GNbp VDD VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=0.36u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=0.36u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=0.36u l=0.1u
mp3 GNb GNbb VDD VDD pmos1v w=0.36u l=0.1u
mp5 n7 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n7 GNbb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATNSRXL

* Spice subcircuit definition for TLATNTSCAX12




.subckt TLATNTSCAX12 ECK / CK E SE
mn0 Eb SE VSS VSS nmos1v w=0.24u l=0.1u
mn1 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n5 VSS VSS nmos1v w=0.43u l=0.1u
mn15 n10 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n10 CKbb n5 VSS nmos1v w=0.24u l=0.1u
mn2 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn20 n15 Eint VSS VSS nmos1v w=1.29u l=0.1u
mn21 n15 CKbb ECKb VSS nmos1v w=1.29u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=5.16u l=0.1u
mn3 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn5 Eb CKb n5 VSS nmos1v w=0.24u l=0.1u
mp0 n0 SE VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 E Eb VDD pmos1v w=0.36u l=0.1u
mp10 Eint n5 VDD VDD pmos1v w=0.65u l=0.1u
mp15 n11 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n11 CKb n5 VDD pmos1v w=0.36u l=0.1u
mp2 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=1.95u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=1.95u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=7.8u l=0.1u
mp3 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp5 Eb CKbb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATNTSCAX12

* Spice subcircuit definition for TLATNTSCAX16




.subckt TLATNTSCAX16 ECK / CK E SE
mn0 Eb SE VSS VSS nmos1v w=0.24u l=0.1u
mn1 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n5 VSS VSS nmos1v w=0.68u l=0.1u
mn15 n10 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n10 CKbb n5 VSS nmos1v w=0.24u l=0.1u
mn2 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn20 n15 Eint VSS VSS nmos1v w=1.72u l=0.1u
mn21 n15 CKbb ECKb VSS nmos1v w=1.72u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=6.88u l=0.1u
mn3 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn5 Eb CKb n5 VSS nmos1v w=0.24u l=0.1u
mp0 n0 SE VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 E Eb VDD pmos1v w=0.36u l=0.1u
mp10 Eint n5 VDD VDD pmos1v w=1.04u l=0.1u
mp15 n11 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n11 CKb n5 VDD pmos1v w=0.36u l=0.1u
mp2 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=2.6u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=2.6u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=10.4u l=0.1u
mp3 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp5 Eb CKbb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATNTSCAX16

* Spice subcircuit definition for TLATNTSCAX2




.subckt TLATNTSCAX2 ECK / CK E SE
mn0 Eb SE VSS VSS nmos1v w=0.24u l=0.1u
mn1 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n5 VSS VSS nmos1v w=0.24u l=0.1u
mn15 n10 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n10 CKbb n5 VSS nmos1v w=0.24u l=0.1u
mn2 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn20 n15 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn21 n15 CKbb ECKb VSS nmos1v w=0.24u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=0.86u l=0.1u
mn3 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn5 Eb CKb n5 VSS nmos1v w=0.24u l=0.1u
mp0 n0 SE VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 E Eb VDD pmos1v w=0.36u l=0.1u
mp10 Eint n5 VDD VDD pmos1v w=0.36u l=0.1u
mp15 n11 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n11 CKb n5 VDD pmos1v w=0.36u l=0.1u
mp2 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=0.36u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=0.36u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=1.3u l=0.1u
mp3 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp5 Eb CKbb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATNTSCAX2

* Spice subcircuit definition for TLATNTSCAX20




.subckt TLATNTSCAX20 ECK / CK E SE
mn0 Eb SE VSS VSS nmos1v w=0.24u l=0.1u
mn1 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n5 VSS VSS nmos1v w=0.86u l=0.1u
mn15 n10 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n10 CKbb n5 VSS nmos1v w=0.24u l=0.1u
mn2 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn20 n15 Eint VSS VSS nmos1v w=2.15u l=0.1u
mn21 n15 CKbb ECKb VSS nmos1v w=2.15u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=8.6u l=0.1u
mn3 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn5 Eb CKb n5 VSS nmos1v w=0.24u l=0.1u
mp0 n0 SE VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 E Eb VDD pmos1v w=0.36u l=0.1u
mp10 Eint n5 VDD VDD pmos1v w=1.3u l=0.1u
mp15 n11 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n11 CKb n5 VDD pmos1v w=0.36u l=0.1u
mp2 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=3.25u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=3.25u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=13.0u l=0.1u
mp3 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp5 Eb CKbb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATNTSCAX20

* Spice subcircuit definition for TLATNTSCAX3




.subckt TLATNTSCAX3 ECK / CK E SE
mn0 Eb SE VSS VSS nmos1v w=0.24u l=0.1u
mn1 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n5 VSS VSS nmos1v w=0.24u l=0.1u
mn15 n10 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n10 CKbb n5 VSS nmos1v w=0.24u l=0.1u
mn2 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn20 n15 Eint VSS VSS nmos1v w=0.43u l=0.1u
mn21 n15 CKbb ECKb VSS nmos1v w=0.43u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=1.29u l=0.1u
mn3 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn5 Eb CKb n5 VSS nmos1v w=0.24u l=0.1u
mp0 n0 SE VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 E Eb VDD pmos1v w=0.36u l=0.1u
mp10 Eint n5 VDD VDD pmos1v w=0.36u l=0.1u
mp15 n11 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n11 CKb n5 VDD pmos1v w=0.36u l=0.1u
mp2 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=0.65u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=0.65u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=1.95u l=0.1u
mp3 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp5 Eb CKbb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATNTSCAX3

* Spice subcircuit definition for TLATNTSCAX4




.subckt TLATNTSCAX4 ECK / CK E SE
mn0 Eb SE VSS VSS nmos1v w=0.24u l=0.1u
mn1 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n5 VSS VSS nmos1v w=0.24u l=0.1u
mn15 n10 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n10 CKbb n5 VSS nmos1v w=0.24u l=0.1u
mn2 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn20 n15 Eint VSS VSS nmos1v w=0.43u l=0.1u
mn21 n15 CKbb ECKb VSS nmos1v w=0.43u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=1.72u l=0.1u
mn3 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn5 Eb CKb n5 VSS nmos1v w=0.24u l=0.1u
mp0 n0 SE VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 E Eb VDD pmos1v w=0.36u l=0.1u
mp10 Eint n5 VDD VDD pmos1v w=0.36u l=0.1u
mp15 n11 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n11 CKb n5 VDD pmos1v w=0.36u l=0.1u
mp2 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=0.65u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=0.65u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=2.6u l=0.1u
mp3 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp5 Eb CKbb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATNTSCAX4

* Spice subcircuit definition for TLATNTSCAX6




.subckt TLATNTSCAX6 ECK / CK E SE
mn0 Eb SE VSS VSS nmos1v w=0.24u l=0.1u
mn1 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n5 VSS VSS nmos1v w=0.34u l=0.1u
mn15 n10 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n10 CKbb n5 VSS nmos1v w=0.24u l=0.1u
mn2 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn20 n15 Eint VSS VSS nmos1v w=0.86u l=0.1u
mn21 n15 CKbb ECKb VSS nmos1v w=0.86u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=2.58u l=0.1u
mn3 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn5 Eb CKb n5 VSS nmos1v w=0.24u l=0.1u
mp0 n0 SE VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 E Eb VDD pmos1v w=0.36u l=0.1u
mp10 Eint n5 VDD VDD pmos1v w=0.52u l=0.1u
mp15 n11 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n11 CKb n5 VDD pmos1v w=0.36u l=0.1u
mp2 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=1.3u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=1.3u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=3.9u l=0.1u
mp3 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp5 Eb CKbb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATNTSCAX6

* Spice subcircuit definition for TLATNTSCAX8




.subckt TLATNTSCAX8 ECK / CK E SE
mn0 Eb SE VSS VSS nmos1v w=0.24u l=0.1u
mn1 Eb E VSS VSS nmos1v w=0.24u l=0.1u
mn10 Eint n5 VSS VSS nmos1v w=0.34u l=0.1u
mn15 n10 Eint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n10 CKbb n5 VSS nmos1v w=0.24u l=0.1u
mn2 CKb CK VSS VSS nmos1v w=0.24u l=0.1u
mn20 n15 Eint VSS VSS nmos1v w=0.86u l=0.1u
mn21 n15 CKbb ECKb VSS nmos1v w=0.86u l=0.1u
mn22 ECK ECKb VSS VSS nmos1v w=3.44u l=0.1u
mn3 CKbb CKb VSS VSS nmos1v w=0.24u l=0.1u
mn5 Eb CKb n5 VSS nmos1v w=0.24u l=0.1u
mp0 n0 SE VDD VDD pmos1v w=0.36u l=0.1u
mp1 n0 E Eb VDD pmos1v w=0.36u l=0.1u
mp10 Eint n5 VDD VDD pmos1v w=0.52u l=0.1u
mp15 n11 Eint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n11 CKb n5 VDD pmos1v w=0.36u l=0.1u
mp2 CKb CK VDD VDD pmos1v w=0.36u l=0.1u
mp20 ECKb Eint VDD VDD pmos1v w=1.3u l=0.1u
mp21 ECKb CKbb VDD VDD pmos1v w=1.3u l=0.1u
mp22 ECK ECKb VDD VDD pmos1v w=5.2u l=0.1u
mp3 CKbb CKb VDD VDD pmos1v w=0.36u l=0.1u
mp5 Eb CKbb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATNTSCAX8

* Spice subcircuit definition for TLATNX1




.subckt TLATNX1 Q QN / D GN
mn0 GNb GN VSS VSS nmos1v w=0.24u l=0.1u
mn1 GNbb GNb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Qint n0 VSS VSS nmos1v w=0.24u l=0.1u
mn15 n5 Qint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 GNbb n0 VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=0.43u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=0.43u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=0.43u l=0.1u
mn5 n1 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 GNb n0 VSS nmos1v w=0.24u l=0.1u
mp0 GNb GN VDD VDD pmos1v w=0.36u l=0.1u
mp1 GNbb GNb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint n0 VDD VDD pmos1v w=0.36u l=0.1u
mp15 n6 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 GNb n0 VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=0.65u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=0.65u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=0.65u l=0.1u
mp5 n2 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 GNbb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATNX1

* Spice subcircuit definition for TLATNX2




.subckt TLATNX2 Q QN / D GN
mn0 GNb GN VSS VSS nmos1v w=0.24u l=0.1u
mn1 GNbb GNb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Qint n0 VSS VSS nmos1v w=0.34u l=0.1u
mn15 n5 Qint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 GNbb n0 VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=0.86u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=0.86u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=0.86u l=0.1u
mn5 n1 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 GNb n0 VSS nmos1v w=0.24u l=0.1u
mp0 GNb GN VDD VDD pmos1v w=0.36u l=0.1u
mp1 GNbb GNb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint n0 VDD VDD pmos1v w=0.52u l=0.1u
mp15 n6 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 GNb n0 VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=1.3u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=1.3u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=1.3u l=0.1u
mp5 n2 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 GNbb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATNX2

* Spice subcircuit definition for TLATNX4




.subckt TLATNX4 Q QN / D GN
mn0 GNb GN VSS VSS nmos1v w=0.24u l=0.1u
mn1 GNbb GNb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Qint n0 VSS VSS nmos1v w=0.68u l=0.1u
mn15 n5 Qint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 GNbb n0 VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=1.72u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=1.72u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=1.72u l=0.1u
mn5 n1 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 GNb n0 VSS nmos1v w=0.24u l=0.1u
mp0 GNb GN VDD VDD pmos1v w=0.36u l=0.1u
mp1 GNbb GNb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint n0 VDD VDD pmos1v w=1.04u l=0.1u
mp15 n6 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 GNb n0 VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=2.6u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=2.6u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=2.6u l=0.1u
mp5 n2 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 GNbb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATNX4

* Spice subcircuit definition for TLATNXL




.subckt TLATNXL Q QN / D GN
mn0 GNb GN VSS VSS nmos1v w=0.24u l=0.1u
mn1 GNbb GNb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Qint n0 VSS VSS nmos1v w=0.24u l=0.1u
mn15 n5 Qint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 GNbb n0 VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=0.24u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=0.24u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=0.24u l=0.1u
mn5 n1 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 GNb n0 VSS nmos1v w=0.24u l=0.1u
mp0 GNb GN VDD VDD pmos1v w=0.36u l=0.1u
mp1 GNbb GNb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint n0 VDD VDD pmos1v w=0.36u l=0.1u
mp15 n6 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 GNb n0 VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=0.36u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=0.36u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=0.36u l=0.1u
mp5 n2 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 GNbb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATNXL

* Spice subcircuit definition for TLATSRX1




.subckt TLATSRX1 Q QN / D G RN SN
mn0 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 G Gb VSS nmos1v w=0.24u l=0.1u
mn10 n10 SN VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 n5 Qint VSS nmos1v w=0.24u l=0.1u
mn15 n17 RN VSS VSS nmos1v w=0.24u l=0.1u
mn16 n17 Qint n15 VSS nmos1v w=0.24u l=0.1u
mn17 n15 Gb n5 VSS nmos1v w=0.24u l=0.1u
mn2 Gbb Gb VSS VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=0.43u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=0.43u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=0.43u l=0.1u
mn5 n6 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n6 Gbb n5 VSS nmos1v w=0.24u l=0.1u
mp0 Gb RN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Gb G VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint SN VDD VDD pmos1v w=0.36u l=0.1u
mp11 Qint n5 VDD VDD pmos1v w=0.36u l=0.1u
mp15 n16 RN VDD VDD pmos1v w=0.36u l=0.1u
mp16 n16 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp17 n16 Gbb n5 VDD pmos1v w=0.36u l=0.1u
mp2 Gbb Gb VDD VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=0.65u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=0.65u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=0.65u l=0.1u
mp5 n7 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n7 Gb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATSRX1

* Spice subcircuit definition for TLATSRX2




.subckt TLATSRX2 Q QN / D G RN SN
mn0 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 G Gb VSS nmos1v w=0.24u l=0.1u
mn10 n10 SN VSS VSS nmos1v w=0.34u l=0.1u
mn11 n10 n5 Qint VSS nmos1v w=0.34u l=0.1u
mn15 n17 RN VSS VSS nmos1v w=0.24u l=0.1u
mn16 n17 Qint n15 VSS nmos1v w=0.24u l=0.1u
mn17 n15 Gb n5 VSS nmos1v w=0.24u l=0.1u
mn2 Gbb Gb VSS VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=0.86u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=0.86u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=0.86u l=0.1u
mn5 n6 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n6 Gbb n5 VSS nmos1v w=0.24u l=0.1u
mp0 Gb RN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Gb G VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint SN VDD VDD pmos1v w=0.52u l=0.1u
mp11 Qint n5 VDD VDD pmos1v w=0.52u l=0.1u
mp15 n16 RN VDD VDD pmos1v w=0.36u l=0.1u
mp16 n16 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp17 n16 Gbb n5 VDD pmos1v w=0.36u l=0.1u
mp2 Gbb Gb VDD VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=1.3u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=1.3u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=1.3u l=0.1u
mp5 n7 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n7 Gb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATSRX2

* Spice subcircuit definition for TLATSRX4




.subckt TLATSRX4 Q QN / D G RN SN
mn0 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 G Gb VSS nmos1v w=0.24u l=0.1u
mn10 n10 SN VSS VSS nmos1v w=0.68u l=0.1u
mn11 n10 n5 Qint VSS nmos1v w=0.68u l=0.1u
mn15 n17 RN VSS VSS nmos1v w=0.24u l=0.1u
mn16 n17 Qint n15 VSS nmos1v w=0.24u l=0.1u
mn17 n15 Gb n5 VSS nmos1v w=0.24u l=0.1u
mn2 Gbb Gb VSS VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=1.72u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=1.72u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=1.72u l=0.1u
mn5 n6 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n6 Gbb n5 VSS nmos1v w=0.24u l=0.1u
mp0 Gb RN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Gb G VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint SN VDD VDD pmos1v w=1.04u l=0.1u
mp11 Qint n5 VDD VDD pmos1v w=1.04u l=0.1u
mp15 n16 RN VDD VDD pmos1v w=0.36u l=0.1u
mp16 n16 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp17 n16 Gbb n5 VDD pmos1v w=0.36u l=0.1u
mp2 Gbb Gb VDD VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=2.6u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=2.6u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=2.6u l=0.1u
mp5 n7 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n7 Gb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATSRX4

* Spice subcircuit definition for TLATSRXL




.subckt TLATSRXL Q QN / D G RN SN
mn0 n0 RN VSS VSS nmos1v w=0.24u l=0.1u
mn1 n0 G Gb VSS nmos1v w=0.24u l=0.1u
mn10 n10 SN VSS VSS nmos1v w=0.24u l=0.1u
mn11 n10 n5 Qint VSS nmos1v w=0.24u l=0.1u
mn15 n17 RN VSS VSS nmos1v w=0.24u l=0.1u
mn16 n17 Qint n15 VSS nmos1v w=0.24u l=0.1u
mn17 n15 Gb n5 VSS nmos1v w=0.24u l=0.1u
mn2 Gbb Gb VSS VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=0.24u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=0.24u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=0.24u l=0.1u
mn5 n6 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n6 Gbb n5 VSS nmos1v w=0.24u l=0.1u
mp0 Gb RN VDD VDD pmos1v w=0.36u l=0.1u
mp1 Gb G VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint SN VDD VDD pmos1v w=0.36u l=0.1u
mp11 Qint n5 VDD VDD pmos1v w=0.36u l=0.1u
mp15 n16 RN VDD VDD pmos1v w=0.36u l=0.1u
mp16 n16 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp17 n16 Gbb n5 VDD pmos1v w=0.36u l=0.1u
mp2 Gbb Gb VDD VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=0.36u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=0.36u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=0.36u l=0.1u
mp5 n7 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n7 Gb n5 VDD pmos1v w=0.36u l=0.1u
.ends TLATSRXL

* Spice subcircuit definition for TLATX1




.subckt TLATX1 Q QN / D G
mn0 Gb G VSS VSS nmos1v w=0.24u l=0.1u
mn1 Gbb Gb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Qint n0 VSS VSS nmos1v w=0.24u l=0.1u
mn15 n5 Qint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 Gb n0 VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=0.43u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=0.43u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=0.43u l=0.1u
mn5 n1 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 Gbb n0 VSS nmos1v w=0.24u l=0.1u
mp0 Gb G VDD VDD pmos1v w=0.36u l=0.1u
mp1 Gbb Gb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint n0 VDD VDD pmos1v w=0.36u l=0.1u
mp15 n6 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 Gbb n0 VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=0.65u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=0.65u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=0.65u l=0.1u
mp5 n2 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 Gb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATX1

* Spice subcircuit definition for TLATX2




.subckt TLATX2 Q QN / D G
mn0 Gb G VSS VSS nmos1v w=0.24u l=0.1u
mn1 Gbb Gb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Qint n0 VSS VSS nmos1v w=0.34u l=0.1u
mn15 n5 Qint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 Gb n0 VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=0.86u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=0.86u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=0.86u l=0.1u
mn5 n1 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 Gbb n0 VSS nmos1v w=0.24u l=0.1u
mp0 Gb G VDD VDD pmos1v w=0.36u l=0.1u
mp1 Gbb Gb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint n0 VDD VDD pmos1v w=0.52u l=0.1u
mp15 n6 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 Gbb n0 VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=1.3u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=1.3u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=1.3u l=0.1u
mp5 n2 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 Gb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATX2

* Spice subcircuit definition for TLATX4




.subckt TLATX4 Q QN / D G
mn0 Gb G VSS VSS nmos1v w=0.24u l=0.1u
mn1 Gbb Gb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Qint n0 VSS VSS nmos1v w=0.68u l=0.1u
mn15 n5 Qint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 Gb n0 VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=1.72u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=1.72u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=1.72u l=0.1u
mn5 n1 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 Gbb n0 VSS nmos1v w=0.24u l=0.1u
mp0 Gb G VDD VDD pmos1v w=0.36u l=0.1u
mp1 Gbb Gb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint n0 VDD VDD pmos1v w=1.04u l=0.1u
mp15 n6 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 Gbb n0 VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=2.6u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=2.6u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=2.6u l=0.1u
mp5 n2 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 Gb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATX4

* Spice subcircuit definition for TLATXL




.subckt TLATXL Q QN / D G
mn0 Gb G VSS VSS nmos1v w=0.24u l=0.1u
mn1 Gbb Gb VSS VSS nmos1v w=0.24u l=0.1u
mn10 Qint n0 VSS VSS nmos1v w=0.24u l=0.1u
mn15 n5 Qint VSS VSS nmos1v w=0.24u l=0.1u
mn16 n5 Gb n0 VSS nmos1v w=0.24u l=0.1u
mn20 Qbint Qint VSS VSS nmos1v w=0.24u l=0.1u
mn21 Q Qbint VSS VSS nmos1v w=0.24u l=0.1u
mn22 QN Qint VSS VSS nmos1v w=0.24u l=0.1u
mn5 n1 D VSS VSS nmos1v w=0.24u l=0.1u
mn6 n1 Gbb n0 VSS nmos1v w=0.24u l=0.1u
mp0 Gb G VDD VDD pmos1v w=0.36u l=0.1u
mp1 Gbb Gb VDD VDD pmos1v w=0.36u l=0.1u
mp10 Qint n0 VDD VDD pmos1v w=0.36u l=0.1u
mp15 n6 Qint VDD VDD pmos1v w=0.36u l=0.1u
mp16 n6 Gbb n0 VDD pmos1v w=0.36u l=0.1u
mp20 Qbint Qint VDD VDD pmos1v w=0.36u l=0.1u
mp21 Q Qbint VDD VDD pmos1v w=0.36u l=0.1u
mp22 QN Qint VDD VDD pmos1v w=0.36u l=0.1u
mp5 n2 D VDD VDD pmos1v w=0.36u l=0.1u
mp6 n2 Gb n0 VDD pmos1v w=0.36u l=0.1u
.ends TLATXL

* Spice subcircuit definition for XNOR2X1




.subckt XNOR2X1 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n2 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 n2 n0 VSS nmos1v w=0.24u l=0.1u
mn4 n1 B n0 VSS nmos1v w=0.24u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 B n0 VDD pmos1v w=0.36u l=0.1u
mp4 n1 n2 n0 VDD pmos1v w=0.36u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends XNOR2X1

* Spice subcircuit definition for XNOR2X2




.subckt XNOR2X2 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n2 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 n2 n0 VSS nmos1v w=0.24u l=0.1u
mn4 n1 B n0 VSS nmos1v w=0.24u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 B n0 VDD pmos1v w=0.36u l=0.1u
mp4 n1 n2 n0 VDD pmos1v w=0.36u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends XNOR2X2

* Spice subcircuit definition for XNOR2X4




.subckt XNOR2X4 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n2 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 n1 VSS VSS nmos1v w=0.43u l=0.1u
mn3 n3 n2 n0 VSS nmos1v w=0.43u l=0.1u
mn4 n1 B n0 VSS nmos1v w=0.43u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 n1 VDD VDD pmos1v w=0.65u l=0.1u
mp3 n4 B n0 VDD pmos1v w=0.65u l=0.1u
mp4 n1 n2 n0 VDD pmos1v w=0.65u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends XNOR2X4

* Spice subcircuit definition for XNOR2XL




.subckt XNOR2XL Y / A B
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n2 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 n2 n0 VSS nmos1v w=0.24u l=0.1u
mn4 n1 B n0 VSS nmos1v w=0.24u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 B n0 VDD pmos1v w=0.36u l=0.1u
mp4 n1 n2 n0 VDD pmos1v w=0.36u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
.ends XNOR2XL

* Spice subcircuit definition for XOR2X1




.subckt XOR2X1 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n2 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 B n0 VSS nmos1v w=0.24u l=0.1u
mn4 n1 n2 n0 VSS nmos1v w=0.24u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=0.43u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 n2 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n1 B n0 VDD pmos1v w=0.36u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=0.65u l=0.1u
.ends XOR2X1

* Spice subcircuit definition for XOR2X2




.subckt XOR2X2 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n2 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 B n0 VSS nmos1v w=0.24u l=0.1u
mn4 n1 n2 n0 VSS nmos1v w=0.24u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=0.86u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 n2 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n1 B n0 VDD pmos1v w=0.36u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=1.3u l=0.1u
.ends XOR2X2

* Spice subcircuit definition for XOR2X4




.subckt XOR2X4 Y / A B
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n2 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 n1 VSS VSS nmos1v w=0.43u l=0.1u
mn3 n3 B n0 VSS nmos1v w=0.43u l=0.1u
mn4 n1 n2 n0 VSS nmos1v w=0.43u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=1.72u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 n1 VDD VDD pmos1v w=0.65u l=0.1u
mp3 n4 n2 n0 VDD pmos1v w=0.65u l=0.1u
mp4 n1 B n0 VDD pmos1v w=0.65u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=2.6u l=0.1u
.ends XOR2X4

* Spice subcircuit definition for XOR2XL




.subckt XOR2XL Y / A B
mn0 n1 A VSS VSS nmos1v w=0.24u l=0.1u
mn1 n2 B VSS VSS nmos1v w=0.24u l=0.1u
mn2 n3 n1 VSS VSS nmos1v w=0.24u l=0.1u
mn3 n3 B n0 VSS nmos1v w=0.24u l=0.1u
mn4 n1 n2 n0 VSS nmos1v w=0.24u l=0.1u
mn5 Y n0 VSS VSS nmos1v w=0.24u l=0.1u
mp0 n1 A VDD VDD pmos1v w=0.36u l=0.1u
mp1 n2 B VDD VDD pmos1v w=0.36u l=0.1u
mp2 n4 n1 VDD VDD pmos1v w=0.36u l=0.1u
mp3 n4 n2 n0 VDD pmos1v w=0.36u l=0.1u
mp4 n1 B n0 VDD pmos1v w=0.36u l=0.1u
mp5 Y n0 VDD VDD pmos1v w=0.36u l=0.1u
.ends XOR2XL

* Spice subcircuit definition for ACHCONX2


.subckt ACHCONX2 CON / A B CI
mn1 n10 n13 n11 VSS nmos1v w=0.52u l=0.1u
mn10 n14 CI VSS VSS nmos1v w=0.65u l=0.1u
mn11 n13 B VSS VSS nmos1v w=0.65u l=0.1u
mn2 n10 B n15 VSS nmos1v w=0.65u l=0.1u
mn3 n9 n13 n15 VSS nmos1v w=0.65u l=0.1u
mn4 n9 B n11 VSS nmos1v w=0.52u l=0.1u
mn5 n11 n15 VSS VSS nmos1v w=0.52u l=0.1u
mn6 n15 A VSS VSS nmos1v w=0.65u l=0.1u
mn7 n12 B VSS VSS nmos1v w=0.65u l=0.1u
mn8 CON n10 n14 VSS nmos1v w=0.65u l=0.1u
mn9 CON n9 n12 VSS nmos1v w=0.65u l=0.1u
mp1 n10 B n11 VDD pmos1v w=0.86u l=0.1u
mp10 n14 CI VDD VDD pmos1v w=1.29u l=0.1u
mp11 n13 B VDD VDD pmos1v w=1.29u l=0.1u
mp2 n10 n13 n15 VDD pmos1v w=1.29u l=0.1u
mp3 n9 B n15 VDD pmos1v w=1.29u l=0.1u
mp4 n9 n13 n11 VDD pmos1v w=0.86u l=0.1u
mp5 n11 n15 VDD VDD pmos1v w=0.86u l=0.1u
mp6 n15 A VDD VDD pmos1v w=1.29u l=0.1u
mp7 n12 B VDD VDD pmos1v w=1.29u l=0.1u
mp8 CON n9 n14 VDD pmos1v w=1.29u l=0.1u
mp9 CON n10 n12 VDD pmos1v w=1.29u l=0.1u
.ENDS ACHCONX2

* Spice subcircuit definition for XNOR3X1


.subckt XNOR3X1 Y / A B C
mn1 n9 B n8 VSS nmos1v w=0.32u l=0.1u
mn10 n12 n61 n8 VSS nmos1v w=0.34u l=0.1u
mn11 n12 B n62 VSS nmos1v w=0.34u l=0.1u
mn2 n9 n61 n62 VSS nmos1v w=0.34u l=0.1u
mn3 n62 A VSS VSS nmos1v w=0.34u l=0.1u
mn4 n61 B VSS VSS nmos1v w=0.32u l=0.1u
mn5 n11 n60 n12 VSS nmos1v w=0.32u l=0.1u
mn6 n11 C n9 VSS nmos1v w=0.32u l=0.1u
mn7 n60 C VSS VSS nmos1v w=0.32u l=0.1u
mn8 Y n11 VSS VSS nmos1v w=0.34u l=0.1u
mn9 n8 n62 VSS VSS nmos1v w=0.32u l=0.1u
mp1 n9 n61 n8 VDD pmos1v w=0.52u l=0.1u
mp10 n12 B n8 VDD pmos1v w=0.52u l=0.1u
mp11 n12 n61 n62 VDD pmos1v w=0.65u l=0.1u
mp2 n9 B n62 VDD pmos1v w=0.65u l=0.1u
mp3 n62 A VDD VDD pmos1v w=0.65u l=0.1u
mp4 n61 B VDD VDD pmos1v w=0.52u l=0.1u
mp5 n11 C n12 VDD pmos1v w=0.52u l=0.1u
mp6 n11 n60 n9 VDD pmos1v w=0.52u l=0.1u
mp7 n60 C VDD VDD pmos1v w=0.52u l=0.1u
mp8 Y n11 VDD VDD pmos1v w=0.65u l=0.1u
mp9 n8 n62 VDD VDD pmos1v w=0.52u l=0.1u
.ENDS XNOR3X1


* Spice subcircuit definition for XNOR3XL


.subckt XNOR3XL Y / A B C
mn0 n12 B n10 VSS nmos1v w=0.32u l=0.1u
mn1 n9 B n8 VSS nmos1v w=0.32u l=0.1u
mn10 n12 n13 n8 VSS nmos1v w=0.34u l=0.1u
mn2 n9 n13 n10 VSS nmos1v w=0.32u l=0.1u
mn3 n10 A VSS VSS nmos1v w=0.34u l=0.1u
mn4 n13 B VSS VSS nmos1v w=0.32u l=0.1u
mn5 n11 n14 n12 VSS nmos1v w=0.32u l=0.1u
mn6 n11 C n9 VSS nmos1v w=0.32u l=0.1u
mn7 n14 C VSS VSS nmos1v w=0.32u l=0.1u
mn8 Y n11 VSS VSS nmos1v w=0.34u l=0.1u
mn9 n8 n10 VSS VSS nmos1v w=0.32u l=0.1u
mp0 n12 n13 n10 VDD pmos1v w=0.52u l=0.1u
mp1 n9 n13 n8 VDD pmos1v w=0.52u l=0.1u
mp10 n12 B n8 VDD pmos1v w=0.52u l=0.1u
mp2 n9 B n10 VDD pmos1v w=0.52u l=0.1u
mp3 n10 A VDD VDD pmos1v w=0.52u l=0.1u
mp4 n13 B VDD VDD pmos1v w=0.52u l=0.1u
mp5 n11 C n12 VDD pmos1v w=0.52u l=0.1u
mp6 n11 n14 n9 VDD pmos1v w=0.52u l=0.1u
mp7 n14 C VDD VDD pmos1v w=0.52u l=0.1u
mp8 Y n11 VDD VDD pmos1v w=0.34u l=0.1u
mp9 n8 n10 VDD VDD pmos1v w=0.52u l=0.1u
.ENDS XNOR3XL

* Spice subcircuit definition for XOR3X1


.subckt XOR3X1 Y / A B C
mn0 n11 n62 VSS VSS nmos1v w=0.32u l=0.1u
mn1 n44 B n62 VSS nmos1v w=0.34u l=0.1u
mn10 n62 A VSS VSS nmos1v w=0.34u l=0.1u
mn2 n44 n61 n11 VSS nmos1v w=0.32u l=0.1u
mn3 n50 n60 n56 VSS nmos1v w=0.32u l=0.1u
mn4 n50 C n44 VSS nmos1v w=0.32u l=0.1u
mn5 n56 n61 n62 VSS nmos1v w=0.34u l=0.1u
mn6 n56 B n11 VSS nmos1v w=0.32u l=0.1u
mn7 Y n50 VSS VSS nmos1v w=0.34u l=0.1u
mn8 n60 C VSS VSS nmos1v w=0.32u l=0.1u
mn9 n61 B VSS VSS nmos1v w=0.32u l=0.1u
mp0 VDD n62 n11 VDD pmos1v w=0.52u l=0.1u
mp1 n44 n61 n62 VDD pmos1v w=0.65u l=0.1u
mp10 VDD A n62 VDD pmos1v w=0.65u l=0.1u
mp2 n44 B n11 VDD pmos1v w=0.52u l=0.1u
mp3 n50 C n56 VDD pmos1v w=0.52u l=0.1u
mp4 n50 n60 n44 VDD pmos1v w=0.52u l=0.1u
mp5 n56 B n62 VDD pmos1v w=0.65u l=0.1u
mp6 n56 n61 n11 VDD pmos1v w=0.52u l=0.1u
mp7 VDD n50 Y VDD pmos1v w=0.65u l=0.1u
mp8 VDD C n60 VDD pmos1v w=0.52u l=0.1u
mp9 VDD B n61 VDD pmos1v w=0.52u l=0.1u
.ENDS XOR3X1

* Spice subcircuit definition for XOR3XL


.subckt XOR3XL Y / A B C
mn0 n11 n19 VSS VSS nmos1v w=0.32u l=0.1u
mn1 n44 B n19 VSS nmos1v w=0.32u l=0.1u
mn10 n19 A VSS VSS nmos1v w=0.32u l=0.1u
mn2 n44 n17 n11 VSS nmos1v w=0.32u l=0.1u
mn3 n50 n30 n56 VSS nmos1v w=0.32u l=0.1u
mn4 n50 C n44 VSS nmos1v w=0.32u l=0.1u
mn5 n56 n17 n19 VSS nmos1v w=0.32u l=0.1u
mn6 n56 B n11 VSS nmos1v w=0.32u l=0.1u
mn7 Y n50 VSS VSS nmos1v w=0.32u l=0.1u
mn8 n30 C VSS VSS nmos1v w=0.32u l=0.1u
mn9 n17 B VSS VSS nmos1v w=0.32u l=0.1u
mp0 VDD n19 n11 VDD pmos1v w=0.52u l=0.1u
mp1 n44 n17 n19 VDD pmos1v w=0.52u l=0.1u
mp10 VDD A n19 VDD pmos1v w=0.52u l=0.1u
mp2 n44 B n11 VDD pmos1v w=0.52u l=0.1u
mp3 n50 C n56 VDD pmos1v w=0.52u l=0.1u
mp4 n50 n30 n44 VDD pmos1v w=0.52u l=0.1u
mp5 n56 B n19 VDD pmos1v w=0.52u l=0.1u
mp6 n56 n17 n11 VDD pmos1v w=0.52u l=0.1u
mp7 VDD n50 Y VDD pmos1v w=0.34u l=0.1u
mp8 VDD C n30 VDD pmos1v w=0.52u l=0.1u
mp9 VDD B n17 VDD pmos1v w=0.52u l=0.1u
.ENDS XOR3XL


.subckt FILL1
.ENDS FILL1

.subckt FILL2
.ENDS FILL2

.subckt FILL4
.ENDS FILL4

.subckt FILL8
.ENDS FILL8

.subckt FILL16
.ENDS FILL16

.subckt FILL32
.ENDS FILL32

.subckt FILL64
.ENDS FILL64

