VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  CAPACITANCE PICOFARADS 1 ;
  DATABASE MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.005 ;
LAYER Oxide
  TYPE MASTERSLICE ;
END Oxide

LAYER Poly
  TYPE MASTERSLICE ;
END Poly

LAYER Nhvt
  TYPE IMPLANT ;
END Nhvt

LAYER Nimp
  TYPE IMPLANT ;
  WIDTH 0.24 ;
  SPACING 0.24 ;
END Nimp

LAYER Phvt
  TYPE IMPLANT ;
END Phvt

LAYER Pimp
  TYPE IMPLANT ;
  WIDTH 0.24 ;
  SPACING 0.24 ;
  SPACING 0 LAYER Nimp ;
END Pimp

LAYER Nzvt
  TYPE IMPLANT ;
  WIDTH 0.7 ;
  SPACING 0.6 ;
END Nzvt

LAYER SiProt
  TYPE IMPLANT ;
  WIDTH 0.44 ;
  SPACING 0.44 ;
END SiProt

LAYER Cont
  TYPE CUT ;
  SPACING 0.14 ;
  SPACING 0.16 ADJACENTCUTS 3 WITHIN 0.17 ;
  WIDTH 0.12 ;
  ENCLOSURE ABOVE 0 0.06 ;
  ANTENNAMODEL OXIDE1 ;
END Cont

LAYER Metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.29 0.29 ;
  WIDTH 0.12 ;
  AREA 0.07 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.559 1.499 2.999 4.499 7.499 
    WIDTH 0 0.12 0.12 0.12 0.12 0.12 0.12 
    WIDTH 0.18 0.12 0.18 0.18 0.18 0.18 0.18 
    WIDTH 1.5 0.18 0.18 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 2 WIDTH 0.4 ;
  MINIMUMCUT 4 WIDTH 1 ;
  MINIMUMCUT 2 WIDTH 2 LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.08 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.3 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
END Metal1

LAYER Via1
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.2 ADJACENTCUTS 3 WITHIN 0.21 ;
  WIDTH 0.14 ;
  ENCLOSURE BELOW 0.005 0.06 ;
  ENCLOSURE ABOVE 0.005 0.06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
END Via1

LAYER Metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.29 0.29 ;
  WIDTH 0.14 ;
  AREA 0.08 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.559 1.499 2.999 4.499 7.499 
    WIDTH 0 0.14 0.14 0.14 0.14 0.14 0.14 
    WIDTH 0.2 0.14 0.2 0.2 0.2 0.2 0.2 
    WIDTH 1.5 0.2 0.2 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 2 WIDTH 0.4 ;
  MINIMUMCUT 4 WIDTH 1 ;
  MINIMUMCUT 2 WIDTH 2 LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.06 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.36 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
END Metal2

LAYER Via2
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.2 ADJACENTCUTS 3 WITHIN 0.21 ;
  WIDTH 0.14 ;
  ENCLOSURE BELOW 0.005 0.06 ;
  ENCLOSURE ABOVE 0.005 0.06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
END Via2

LAYER Metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.29 0.29 ;
  WIDTH 0.14 ;
  AREA 0.08 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.559 1.499 2.999 4.499 7.499 
    WIDTH 0 0.14 0.14 0.14 0.14 0.14 0.14 
    WIDTH 0.2 0.14 0.2 0.2 0.2 0.2 0.2 
    WIDTH 1.5 0.2 0.2 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 2 WIDTH 0.4 ;
  MINIMUMCUT 4 WIDTH 1 ;
  MINIMUMCUT 2 WIDTH 2 LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.06 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.36 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
END Metal3

LAYER Via3
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.2 ADJACENTCUTS 3 WITHIN 0.21 ;
  WIDTH 0.14 ;
  ENCLOSURE BELOW 0.005 0.06 ;
  ENCLOSURE ABOVE 0.005 0.06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
END Via3

LAYER Metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.29 0.29 ;
  WIDTH 0.14 ;
  AREA 0.08 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.559 1.499 2.999 4.499 7.499 
    WIDTH 0 0.14 0.14 0.14 0.14 0.14 0.14 
    WIDTH 0.2 0.14 0.2 0.2 0.2 0.2 0.2 
    WIDTH 1.5 0.2 0.2 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 2 WIDTH 0.4 ;
  MINIMUMCUT 4 WIDTH 1 ;
  MINIMUMCUT 2 WIDTH 2 LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.06 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.36 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
END Metal4

LAYER Via4
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.2 ADJACENTCUTS 3 WITHIN 0.21 ;
  WIDTH 0.14 ;
  ENCLOSURE BELOW 0.005 0.06 ;
  ENCLOSURE ABOVE 0.005 0.06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
END Via4

LAYER Metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.29 0.29 ;
  WIDTH 0.14 ;
  AREA 0.08 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.559 1.499 2.999 4.499 7.499 
    WIDTH 0 0.14 0.14 0.14 0.14 0.14 0.14 
    WIDTH 0.2 0.14 0.2 0.2 0.2 0.2 0.2 
    WIDTH 1.5 0.2 0.2 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 2 WIDTH 0.4 ;
  MINIMUMCUT 4 WIDTH 1 ;
  MINIMUMCUT 2 WIDTH 2 LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.06 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.36 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
END Metal5

LAYER Via5
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.2 ADJACENTCUTS 3 WITHIN 0.21 ;
  WIDTH 0.14 ;
  ENCLOSURE BELOW 0.005 0.06 ;
  ENCLOSURE ABOVE 0.005 0.06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
END Via5

LAYER Metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.29 0.29 ;
  WIDTH 0.14 ;
  AREA 0.08 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.559 1.499 2.999 4.499 7.499 
    WIDTH 0 0.14 0.14 0.14 0.14 0.14 0.14 
    WIDTH 0.2 0.14 0.2 0.2 0.2 0.2 0.2 
    WIDTH 1.5 0.2 0.2 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 2 WIDTH 0.4 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 1 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 1.6 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 4 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 2 LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.06 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.36 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
END Metal6

LAYER Via6
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.2 ADJACENTCUTS 3 WITHIN 0.21 ;
  WIDTH 0.14 ;
  ENCLOSURE BELOW 0.005 0.06 ;
  ENCLOSURE ABOVE 0.005 0.06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
END Via6

LAYER Metal7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.29 0.29 ;
  WIDTH 0.14 ;
  AREA 0.08 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.559 1.499 2.999 4.499 7.499 
    WIDTH 0 0.14 0.14 0.14 0.14 0.14 0.14 
    WIDTH 0.2 0.14 0.2 0.2 0.2 0.2 0.2 
    WIDTH 1.5 0.2 0.2 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 2 WIDTH 1.6 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 4 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 2 LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.06 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.36 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
END Metal7

LAYER Via7
  TYPE CUT ;
  SPACING 0.36 ;
  SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.55 ;
  WIDTH 0.36 ;
  ENCLOSURE BELOW 0.03 0.08 ;
  ENCLOSURE ABOVE 0.05 0.1 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
END Via7

LAYER Metal8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.87 0.87 ;
  WIDTH 0.44 ;
  AREA 0.2 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 1.499 2.999 4.499 7.499 
    WIDTH 0 0.4 0.4 0.4 0.4 0.4 
    WIDTH 1.5 0.4 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 2 WIDTH 2 LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.02 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 1 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
END Metal8

LAYER Via8
  TYPE CUT ;
  SPACING 0.36 ;
  SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.55 ;
  WIDTH 0.36 ;
  ENCLOSURE BELOW 0.03 0.08 ;
  ENCLOSURE ABOVE 0.05 0.1 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
END Via8

LAYER Metal9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.87 0.87 ;
  WIDTH 0.44 ;
  AREA 0.2 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 1.499 2.999 4.499 7.499 
    WIDTH 0 0.4 0.4 0.4 0.4 0.4 
    WIDTH 1.5 0.4 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.02 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 1 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
END Metal9

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

MAXVIASTACK 4 RANGE Metal1 Metal7 ;
VIARULE M9_M8v GENERATE
  LAYER Metal8 ;
    ENCLOSURE 0.03 0.08 ;
  LAYER Metal9 ;
    ENCLOSURE 0.05 0.1 ;
  LAYER Via8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.72 BY 0.72 ;
END M9_M8v

VIARULE M8_M7v GENERATE
  LAYER Metal7 ;
    ENCLOSURE 0.03 0.08 ;
  LAYER Metal8 ;
    ENCLOSURE 0.05 0.1 ;
  LAYER Via7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.72 BY 0.72 ;
END M8_M7v

VIARULE M7_M6v GENERATE
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal7 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.29 BY 0.29 ;
END M7_M6v

VIARULE M6_M5v GENERATE
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.29 BY 0.29 ;
END M6_M5v

VIARULE M5_M4v GENERATE
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.29 BY 0.29 ;
END M5_M4v

VIARULE M4_M3v GENERATE
  LAYER Metal3 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.29 BY 0.29 ;
END M4_M3v

VIARULE M3_M2v GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal3 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.29 BY 0.29 ;
END M3_M2v

VIARULE M2_M1v GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal2 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.29 BY 0.29 ;
END M2_M1v

VIARULE M1_POv GENERATE
  LAYER Poly ;
    ENCLOSURE 0.04 0.06 ;
  LAYER Metal1 ;
    ENCLOSURE 0 0.06 ;
  LAYER Cont ;
    RECT -0.06 -0.06 0.06 0.06 ;
    SPACING 0.26 BY 0.26 ;
END M1_POv

VIARULE M9_M8 GENERATE
  LAYER Metal8 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER Metal9 ;
    ENCLOSURE 0.1 0.1 ;
  LAYER Via8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.72 BY 0.72 ;
END M9_M8

VIARULE M8_M7 GENERATE
  LAYER Metal7 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER Metal8 ;
    ENCLOSURE 0.1 0.1 ;
  LAYER Via7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.72 BY 0.72 ;
END M8_M7

VIARULE M7_M6 GENERATE
  LAYER Metal6 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Metal7 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M7_M6

VIARULE M6_M5 GENERATE
  LAYER Metal5 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Metal6 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M6_M5

VIARULE M5_M4 GENERATE
  LAYER Metal4 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Metal5 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M5_M4

VIARULE M4_M3 GENERATE
  LAYER Metal3 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Metal4 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M4_M3

VIARULE M3_M2 GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Metal3 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M3_M2

VIARULE M2_M1 GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Metal2 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Via1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M2_M1

VIARULE M1_PO GENERATE
  LAYER Poly ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Metal1 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Cont ;
    RECT -0.06 -0.06 0.06 0.06 ;
    SPACING 0.28 BY 0.28 ;
END M1_PO

VIARULE M9_M8c GENERATE
  LAYER Metal8 ;
    ENCLOSURE 0.03 0.08 ;
  LAYER Metal9 ;
    ENCLOSURE 0.05 0.1 ;
  LAYER Via8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.72 BY 0.72 ;
END M9_M8c

VIARULE M8_M7c GENERATE
  LAYER Metal7 ;
    ENCLOSURE 0.03 0.08 ;
  LAYER Metal8 ;
    ENCLOSURE 0.05 0.1 ;
  LAYER Via7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.72 BY 0.72 ;
END M8_M7c

VIARULE M7_M6c GENERATE
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal7 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M7_M6c

VIARULE M6_M5c GENERATE
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M6_M5c

VIARULE M5_M4c GENERATE
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M5_M4c

VIARULE M4_M3c GENERATE
  LAYER Metal3 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M4_M3c

VIARULE M3_M2c GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal3 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M3_M2c

VIARULE M2_M1c GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal2 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M2_M1c

VIARULE M1_POLYc GENERATE
  LAYER Poly ;
    ENCLOSURE 0.04 0.06 ;
  LAYER Metal1 ;
    ENCLOSURE 0 0.06 ;
  LAYER Cont ;
    RECT -0.06 -0.06 0.06 0.06 ;
    SPACING 0.28 BY 0.28 ;
END M1_POLYc

SPACING
  SAMENET Poly Poly 0.12 ;
  SAMENET Cont Cont 0.14 ;
  SAMENET Metal1 Metal1 0.12 ;
  SAMENET Via1 Via1 0.15 ;
  SAMENET Metal2 Metal2 0.14 ;
  SAMENET Via2 Via2 0.15 ;
  SAMENET Metal3 Metal3 0.14 ;
  SAMENET Via3 Via3 0.15 ;
  SAMENET Metal4 Metal4 0.14 ;
  SAMENET Via4 Via4 0.15 ;
  SAMENET Metal5 Metal5 0.14 ;
  SAMENET Via5 Via5 0.15 ;
  SAMENET Metal6 Metal6 0.14 ;
  SAMENET Via6 Via6 0.15 ;
  SAMENET Metal7 Metal7 0.14 ;
  SAMENET Via7 Via7 0.36 ;
  SAMENET Metal8 Metal8 0.4 ;
  SAMENET Via8 Via8 0.36 ;
  SAMENET Metal9 Metal9 0.4 ;
END SPACING

END LIBRARY
